/*
MIT License

Copyright Anton Oreskin | https://gosudev.de


Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all
copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
SOFTWARE.
*/
module vulkan

pub fn make_api_version(variant u32, major u32, minor u32, patch u32) u32 {
	return (variant << 29) | (major << 22) | (minor << 12) | patch
}

pub const api_version = make_api_version(0, 1, 0, 0) // patch version should always be set to 0
pub const header_version = 330
pub const header_version_complete = make_api_version(0, 1, 4, header_version)

pub fn make_version(major u32, minor u32, patch u32) u32 {
	return (major << 22) | (minor << 12) | patch
}

pub fn version_major(version u32) u32 {
	return version >> 22
}

pub fn version_minor(version u32) u32 {
	return (version >> 12) & 0xFFF
}

pub fn version_patch(version u32) u32 {
	return version & 0xFFF
}

pub fn version_variant(version u32) u32 {
	return version >> 29
}

pub fn api_version_major(version u32) u32 {
	return (version >> 22) & u32(0x7F)
}

pub fn api_version_minor(version u32) u32 {
	return (version >> 12) & u32(0x3FF)
}

pub fn api_version_patch(version u32) u32 {
	return version & u32(0xFFF)
}

pub const api_version_1_0 = make_api_version(0, 1, 0, 0) // patch version should always be set to 0

pub type Bool32 = u32
pub type DeviceAddress = u64
pub type DeviceSize = u64
pub type Flags = u32
pub type SampleMask = u32

// Pointer to VkBuffer_T
pub type Buffer = voidptr

// Pointer to VkImage_T
pub type Image = voidptr

// Pointer to VkInstance_T
pub type Instance = voidptr

// Pointer to VkPhysicalDevice_T
pub type PhysicalDevice = voidptr

// Pointer to VkDevice_T
pub type Device = voidptr

// Pointer to VkQueue_T
pub type Queue = voidptr

// Pointer to VkSemaphore_T
pub type Semaphore = voidptr

// Pointer to VkCommandBuffer_T
pub type CommandBuffer = voidptr

// Pointer to VkFence_T
pub type Fence = voidptr

// Pointer to VkDeviceMemory_T
pub type DeviceMemory = voidptr

// Pointer to VkQueryPool_T
pub type QueryPool = voidptr

// Pointer to VkImageView_T
pub type ImageView = voidptr

// Pointer to VkCommandPool_T
pub type CommandPool = voidptr

// Pointer to VkRenderPass_T
pub type RenderPass = voidptr

// Pointer to VkFramebuffer_T
pub type Framebuffer = voidptr

// Pointer to VkEvent_T
pub type Event = voidptr

// Pointer to VkBufferView_T
pub type BufferView = voidptr

// Pointer to VkShaderModule_T
pub type ShaderModule = voidptr

// Pointer to VkPipelineCache_T
pub type PipelineCache = voidptr

// Pointer to VkPipelineLayout_T
pub type PipelineLayout = voidptr

// Pointer to VkPipeline_T
pub type Pipeline = voidptr

// Pointer to VkDescriptorSetLayout_T
pub type DescriptorSetLayout = voidptr

// Pointer to VkSampler_T
pub type Sampler = voidptr

// Pointer to VkDescriptorSet_T
pub type DescriptorSet = voidptr

// Pointer to VkDescriptorPool_T
pub type DescriptorPool = voidptr

pub const _false = u32(0)
pub const lod_clamp_none = f32(1000.0)
pub const queue_family_ignored = ~u32(0)
pub const remaining_array_layers = ~u32(0)
pub const remaining_mip_levels = ~u32(0)
pub const _true = u32(1)
pub const whole_size = ~u64(0)
pub const max_memory_types = u32(32)
pub const max_physical_device_name_size = u32(256)
pub const uuid_size = u32(16)
pub const max_extension_name_size = u32(256)
pub const max_description_size = u32(256)
pub const max_memory_heaps = u32(16)
pub const attachment_unused = ~u32(0)
pub const subpass_external = ~u32(0)

pub enum Result {
	success                                            = 0
	not_ready                                          = 1
	timeout                                            = 2
	event_set                                          = 3
	event_reset                                        = 4
	incomplete                                         = 5
	error_out_of_host_memory                           = -1
	error_out_of_device_memory                         = -2
	error_initialization_failed                        = -3
	error_device_lost                                  = -4
	error_memory_map_failed                            = -5
	error_layer_not_present                            = -6
	error_extension_not_present                        = -7
	error_feature_not_present                          = -8
	error_incompatible_driver                          = -9
	error_too_many_objects                             = -10
	error_format_not_supported                         = -11
	error_fragmented_pool                              = -12
	error_unknown                                      = -13
	error_validation_failed                            = -1000011001
	error_out_of_pool_memory                           = -1000069000
	error_invalid_external_handle                      = -1000072003
	error_invalid_opaque_capture_address               = -1000257000
	error_fragmentation                                = -1000161000
	pipeline_compile_required                          = 1000297000
	error_not_permitted                                = -1000174001
	error_surface_lost_khr                             = -1000000000
	error_native_window_in_use_khr                     = -1000000001
	suboptimal_khr                                     = 1000001003
	error_out_of_date_khr                              = -1000001004
	error_incompatible_display_khr                     = -1000003001
	error_invalid_shader_nv                            = -1000012000
	error_image_usage_not_supported_khr                = -1000023000
	error_video_picture_layout_not_supported_khr       = -1000023001
	error_video_profile_operation_not_supported_khr    = -1000023002
	error_video_profile_format_not_supported_khr       = -1000023003
	error_video_profile_codec_not_supported_khr        = -1000023004
	error_video_std_version_not_supported_khr          = -1000023005
	error_invalid_drm_format_modifier_plane_layout_ext = -1000158000
	error_full_screen_exclusive_mode_lost_ext          = -1000255000
	thread_idle_khr                                    = 1000268000
	thread_done_khr                                    = 1000268001
	operation_deferred_khr                             = 1000268002
	operation_not_deferred_khr                         = 1000268003
	error_invalid_video_std_parameters_khr             = -1000299000
	error_compression_exhausted_ext                    = -1000338000
	incompatible_shader_binary_ext                     = 1000482000
	pipeline_binary_missing_khr                        = 1000483000
	error_not_enough_space_khr                         = -1000483000
	max_enum                                           = max_int
}

pub enum StructureType as u32 {
	application_info                                                      = 0
	instance_create_info                                                  = 1
	device_queue_create_info                                              = 2
	device_create_info                                                    = 3
	submit_info                                                           = 4
	memory_allocate_info                                                  = 5
	mapped_memory_range                                                   = 6
	bind_sparse_info                                                      = 7
	fence_create_info                                                     = 8
	semaphore_create_info                                                 = 9
	event_create_info                                                     = 10
	query_pool_create_info                                                = 11
	buffer_create_info                                                    = 12
	buffer_view_create_info                                               = 13
	image_create_info                                                     = 14
	image_view_create_info                                                = 15
	shader_module_create_info                                             = 16
	pipeline_cache_create_info                                            = 17
	pipeline_shader_stage_create_info                                     = 18
	pipeline_vertex_input_state_create_info                               = 19
	pipeline_input_assembly_state_create_info                             = 20
	pipeline_tessellation_state_create_info                               = 21
	pipeline_viewport_state_create_info                                   = 22
	pipeline_rasterization_state_create_info                              = 23
	pipeline_multisample_state_create_info                                = 24
	pipeline_depth_stencil_state_create_info                              = 25
	pipeline_color_blend_state_create_info                                = 26
	pipeline_dynamic_state_create_info                                    = 27
	graphics_pipeline_create_info                                         = 28
	compute_pipeline_create_info                                          = 29
	pipeline_layout_create_info                                           = 30
	sampler_create_info                                                   = 31
	descriptor_set_layout_create_info                                     = 32
	descriptor_pool_create_info                                           = 33
	descriptor_set_allocate_info                                          = 34
	write_descriptor_set                                                  = 35
	copy_descriptor_set                                                   = 36
	framebuffer_create_info                                               = 37
	render_pass_create_info                                               = 38
	command_pool_create_info                                              = 39
	command_buffer_allocate_info                                          = 40
	command_buffer_inheritance_info                                       = 41
	command_buffer_begin_info                                             = 42
	render_pass_begin_info                                                = 43
	buffer_memory_barrier                                                 = 44
	image_memory_barrier                                                  = 45
	memory_barrier                                                        = 46
	loader_instance_create_info                                           = 47
	loader_device_create_info                                             = 48
	bind_buffer_memory_info                                               = 1000157000
	bind_image_memory_info                                                = 1000157001
	memory_dedicated_requirements                                         = 1000127000
	memory_dedicated_allocate_info                                        = 1000127001
	memory_allocate_flags_info                                            = 1000060000
	device_group_command_buffer_begin_info                                = 1000060004
	device_group_submit_info                                              = 1000060005
	device_group_bind_sparse_info                                         = 1000060006
	bind_buffer_memory_device_group_info                                  = 1000060013
	bind_image_memory_device_group_info                                   = 1000060014
	physical_device_group_properties                                      = 1000070000
	device_group_device_create_info                                       = 1000070001
	buffer_memory_requirements_info2                                      = 1000146000
	image_memory_requirements_info2                                       = 1000146001
	image_sparse_memory_requirements_info2                                = 1000146002
	memory_requirements2                                                  = 1000146003
	sparse_image_memory_requirements2                                     = 1000146004
	physical_device_features2                                             = 1000059000
	physical_device_properties2                                           = 1000059001
	format_properties2                                                    = 1000059002
	image_format_properties2                                              = 1000059003
	physical_device_image_format_info2                                    = 1000059004
	queue_family_properties2                                              = 1000059005
	physical_device_memory_properties2                                    = 1000059006
	sparse_image_format_properties2                                       = 1000059007
	physical_device_sparse_image_format_info2                             = 1000059008
	image_view_usage_create_info                                          = 1000117002
	protected_submit_info                                                 = 1000145000
	physical_device_protected_memory_features                             = 1000145001
	physical_device_protected_memory_properties                           = 1000145002
	device_queue_info2                                                    = 1000145003
	physical_device_external_image_format_info                            = 1000071000
	external_image_format_properties                                      = 1000071001
	physical_device_external_buffer_info                                  = 1000071002
	external_buffer_properties                                            = 1000071003
	physical_device_id_properties                                         = 1000071004
	external_memory_buffer_create_info                                    = 1000072000
	external_memory_image_create_info                                     = 1000072001
	export_memory_allocate_info                                           = 1000072002
	physical_device_external_fence_info                                   = 1000112000
	external_fence_properties                                             = 1000112001
	export_fence_create_info                                              = 1000113000
	export_semaphore_create_info                                          = 1000077000
	physical_device_external_semaphore_info                               = 1000076000
	external_semaphore_properties                                         = 1000076001
	physical_device_subgroup_properties                                   = 1000094000
	physical_device16bit_storage_features                                 = 1000083000
	physical_device_variable_pointers_features                            = 1000120000
	descriptor_update_template_create_info                                = 1000085000
	physical_device_maintenance3_properties                               = 1000168000
	descriptor_set_layout_support                                         = 1000168001
	sampler_ycbcr_conversion_create_info                                  = 1000156000
	sampler_ycbcr_conversion_info                                         = 1000156001
	bind_image_plane_memory_info                                          = 1000156002
	image_plane_memory_requirements_info                                  = 1000156003
	physical_device_sampler_ycbcr_conversion_features                     = 1000156004
	sampler_ycbcr_conversion_image_format_properties                      = 1000156005
	device_group_render_pass_begin_info                                   = 1000060003
	physical_device_point_clipping_properties                             = 1000117000
	render_pass_input_attachment_aspect_create_info                       = 1000117001
	pipeline_tessellation_domain_origin_state_create_info                 = 1000117003
	render_pass_multiview_create_info                                     = 1000053000
	physical_device_multiview_features                                    = 1000053001
	physical_device_multiview_properties                                  = 1000053002
	physical_device_shader_draw_parameters_features                       = 1000063000
	physical_device_vulkan1_1_features                                    = 49
	physical_device_vulkan1_1_properties                                  = 50
	physical_device_vulkan1_2_features                                    = 51
	physical_device_vulkan1_2_properties                                  = 52
	image_format_list_create_info                                         = 1000147000
	physical_device_driver_properties                                     = 1000196000
	physical_device_vulkan_memory_model_features                          = 1000211000
	physical_device_host_query_reset_features                             = 1000261000
	physical_device_timeline_semaphore_features                           = 1000207000
	physical_device_timeline_semaphore_properties                         = 1000207001
	semaphore_type_create_info                                            = 1000207002
	timeline_semaphore_submit_info                                        = 1000207003
	semaphore_wait_info                                                   = 1000207004
	semaphore_signal_info                                                 = 1000207005
	physical_device_buffer_device_address_features                        = 1000257000
	buffer_device_address_info                                            = 1000244001
	buffer_opaque_capture_address_create_info                             = 1000257002
	memory_opaque_capture_address_allocate_info                           = 1000257003
	device_memory_opaque_capture_address_info                             = 1000257004
	physical_device8bit_storage_features                                  = 1000177000
	physical_device_shader_atomic_int64_features                          = 1000180000
	physical_device_shader_float16_int8_features                          = 1000082000
	physical_device_float_controls_properties                             = 1000197000
	descriptor_set_layout_binding_flags_create_info                       = 1000161000
	physical_device_descriptor_indexing_features                          = 1000161001
	physical_device_descriptor_indexing_properties                        = 1000161002
	descriptor_set_variable_descriptor_count_allocate_info                = 1000161003
	descriptor_set_variable_descriptor_count_layout_support               = 1000161004
	physical_device_scalar_block_layout_features                          = 1000221000
	physical_device_sampler_filter_minmax_properties                      = 1000130000
	sampler_reduction_mode_create_info                                    = 1000130001
	physical_device_uniform_buffer_standard_layout_features               = 1000253000
	physical_device_shader_subgroup_extended_types_features               = 1000175000
	attachment_description2                                               = 1000109000
	attachment_reference2                                                 = 1000109001
	subpass_description2                                                  = 1000109002
	subpass_dependency2                                                   = 1000109003
	render_pass_create_info2                                              = 1000109004
	subpass_begin_info                                                    = 1000109005
	subpass_end_info                                                      = 1000109006
	physical_device_depth_stencil_resolve_properties                      = 1000199000
	subpass_description_depth_stencil_resolve                             = 1000199001
	image_stencil_usage_create_info                                       = 1000246000
	physical_device_imageless_framebuffer_features                        = 1000108000
	framebuffer_attachments_create_info                                   = 1000108001
	framebuffer_attachment_image_info                                     = 1000108002
	render_pass_attachment_begin_info                                     = 1000108003
	physical_device_separate_depth_stencil_layouts_features               = 1000241000
	attachment_reference_stencil_layout                                   = 1000241001
	attachment_description_stencil_layout                                 = 1000241002
	physical_device_vulkan1_3_features                                    = 53
	physical_device_vulkan1_3_properties                                  = 54
	physical_device_tool_properties                                       = 1000245000
	physical_device_private_data_features                                 = 1000295000
	device_private_data_create_info                                       = 1000295001
	private_data_slot_create_info                                         = 1000295002
	memory_barrier2                                                       = 1000314000
	buffer_memory_barrier2                                                = 1000314001
	image_memory_barrier2                                                 = 1000314002
	dependency_info                                                       = 1000314003
	submit_info2                                                          = 1000314004
	semaphore_submit_info                                                 = 1000314005
	command_buffer_submit_info                                            = 1000314006
	physical_device_synchronization2_features                             = 1000314007
	copy_buffer_info2                                                     = 1000337000
	copy_image_info2                                                      = 1000337001
	copy_buffer_to_image_info2                                            = 1000337002
	copy_image_to_buffer_info2                                            = 1000337003
	buffer_copy2                                                          = 1000337006
	image_copy2                                                           = 1000337007
	buffer_image_copy2                                                    = 1000337009
	physical_device_texture_compression_astc_hdr_features                 = 1000066000
	format_properties3                                                    = 1000360000
	physical_device_maintenance4_features                                 = 1000413000
	physical_device_maintenance4_properties                               = 1000413001
	device_buffer_memory_requirements                                     = 1000413002
	device_image_memory_requirements                                      = 1000413003
	pipeline_creation_feedback_create_info                                = 1000192000
	physical_device_shader_terminate_invocation_features                  = 1000215000
	physical_device_shader_demote_to_helper_invocation_features           = 1000276000
	physical_device_pipeline_creation_cache_control_features              = 1000297000
	physical_device_zero_initialize_workgroup_memory_features             = 1000325000
	physical_device_image_robustness_features                             = 1000335000
	physical_device_subgroup_size_control_properties                      = 1000225000
	pipeline_shader_stage_required_subgroup_size_create_info              = 1000225001
	physical_device_subgroup_size_control_features                        = 1000225002
	physical_device_inline_uniform_block_features                         = 1000138000
	physical_device_inline_uniform_block_properties                       = 1000138001
	write_descriptor_set_inline_uniform_block                             = 1000138002
	descriptor_pool_inline_uniform_block_create_info                      = 1000138003
	physical_device_shader_integer_dot_product_features                   = 1000280000
	physical_device_shader_integer_dot_product_properties                 = 1000280001
	physical_device_texel_buffer_alignment_properties                     = 1000281001
	blit_image_info2                                                      = 1000337004
	resolve_image_info2                                                   = 1000337005
	image_blit2                                                           = 1000337008
	image_resolve2                                                        = 1000337010
	rendering_info                                                        = 1000044000
	rendering_attachment_info                                             = 1000044001
	pipeline_rendering_create_info                                        = 1000044002
	physical_device_dynamic_rendering_features                            = 1000044003
	command_buffer_inheritance_rendering_info                             = 1000044004
	physical_device_vulkan1_4_features                                    = 55
	physical_device_vulkan1_4_properties                                  = 56
	device_queue_global_priority_create_info                              = 1000174000
	physical_device_global_priority_query_features                        = 1000388000
	queue_family_global_priority_properties                               = 1000388001
	physical_device_index_type_uint8_features                             = 1000265000
	memory_map_info                                                       = 1000271000
	memory_unmap_info                                                     = 1000271001
	physical_device_maintenance5_features                                 = 1000470000
	physical_device_maintenance5_properties                               = 1000470001
	device_image_subresource_info                                         = 1000470004
	subresource_layout2                                                   = 1000338002
	image_subresource2                                                    = 1000338003
	buffer_usage_flags2_create_info                                       = 1000470006
	physical_device_maintenance6_features                                 = 1000545000
	physical_device_maintenance6_properties                               = 1000545001
	bind_memory_status                                                    = 1000545002
	physical_device_host_image_copy_features                              = 1000270000
	physical_device_host_image_copy_properties                            = 1000270001
	memory_to_image_copy                                                  = 1000270002
	image_to_memory_copy                                                  = 1000270003
	copy_image_to_memory_info                                             = 1000270004
	copy_memory_to_image_info                                             = 1000270005
	host_image_layout_transition_info                                     = 1000270006
	copy_image_to_image_info                                              = 1000270007
	subresource_host_memcpy_size                                          = 1000270008
	host_image_copy_device_performance_query                              = 1000270009
	physical_device_shader_subgroup_rotate_features                       = 1000416000
	physical_device_shader_float_controls2_features                       = 1000528000
	physical_device_shader_expect_assume_features                         = 1000544000
	pipeline_create_flags2_create_info                                    = 1000470005
	physical_device_push_descriptor_properties                            = 1000080000
	bind_descriptor_sets_info                                             = 1000545003
	push_constants_info                                                   = 1000545004
	push_descriptor_set_info                                              = 1000545005
	push_descriptor_set_with_template_info                                = 1000545006
	physical_device_pipeline_protected_access_features                    = 1000466000
	pipeline_robustness_create_info                                       = 1000068000
	physical_device_pipeline_robustness_features                          = 1000068001
	physical_device_pipeline_robustness_properties                        = 1000068002
	physical_device_line_rasterization_features                           = 1000259000
	pipeline_rasterization_line_state_create_info                         = 1000259001
	physical_device_line_rasterization_properties                         = 1000259002
	physical_device_vertex_attribute_divisor_properties                   = 1000525000
	pipeline_vertex_input_divisor_state_create_info                       = 1000190001
	physical_device_vertex_attribute_divisor_features                     = 1000190002
	rendering_area_info                                                   = 1000470003
	physical_device_dynamic_rendering_local_read_features                 = 1000232000
	rendering_attachment_location_info                                    = 1000232001
	rendering_input_attachment_index_info                                 = 1000232002
	swapchain_create_info_khr                                             = 1000001000
	present_info_khr                                                      = 1000001001
	device_group_present_capabilities_khr                                 = 1000060007
	image_swapchain_create_info_khr                                       = 1000060008
	bind_image_memory_swapchain_info_khr                                  = 1000060009
	acquire_next_image_info_khr                                           = 1000060010
	device_group_present_info_khr                                         = 1000060011
	device_group_swapchain_create_info_khr                                = 1000060012
	display_mode_create_info_khr                                          = 1000002000
	display_surface_create_info_khr                                       = 1000002001
	display_present_info_khr                                              = 1000003000
	xlib_surface_create_info_khr                                          = 1000004000
	xcb_surface_create_info_khr                                           = 1000005000
	wayland_surface_create_info_khr                                       = 1000006000
	android_surface_create_info_khr                                       = 1000008000
	win32_surface_create_info_khr                                         = 1000009000
	debug_report_callback_create_info_ext                                 = 1000011000
	pipeline_rasterization_state_rasterization_order_amd                  = 1000018000
	debug_marker_object_name_info_ext                                     = 1000022000
	debug_marker_object_tag_info_ext                                      = 1000022001
	debug_marker_marker_info_ext                                          = 1000022002
	video_profile_info_khr                                                = 1000023000
	video_capabilities_khr                                                = 1000023001
	video_picture_resource_info_khr                                       = 1000023002
	video_session_memory_requirements_khr                                 = 1000023003
	bind_video_session_memory_info_khr                                    = 1000023004
	video_session_create_info_khr                                         = 1000023005
	video_session_parameters_create_info_khr                              = 1000023006
	video_session_parameters_update_info_khr                              = 1000023007
	video_begin_coding_info_khr                                           = 1000023008
	video_end_coding_info_khr                                             = 1000023009
	video_coding_control_info_khr                                         = 1000023010
	video_reference_slot_info_khr                                         = 1000023011
	queue_family_video_properties_khr                                     = 1000023012
	video_profile_list_info_khr                                           = 1000023013
	physical_device_video_format_info_khr                                 = 1000023014
	video_format_properties_khr                                           = 1000023015
	queue_family_query_result_status_properties_khr                       = 1000023016
	video_decode_info_khr                                                 = 1000024000
	video_decode_capabilities_khr                                         = 1000024001
	video_decode_usage_info_khr                                           = 1000024002
	dedicated_allocation_image_create_info_nv                             = 1000026000
	dedicated_allocation_buffer_create_info_nv                            = 1000026001
	dedicated_allocation_memory_allocate_info_nv                          = 1000026002
	physical_device_transform_feedback_features_ext                       = 1000028000
	physical_device_transform_feedback_properties_ext                     = 1000028001
	pipeline_rasterization_state_stream_create_info_ext                   = 1000028002
	cu_module_create_info_nvx                                             = 1000029000
	cu_function_create_info_nvx                                           = 1000029001
	cu_launch_info_nvx                                                    = 1000029002
	cu_module_texturing_mode_create_info_nvx                              = 1000029004
	image_view_handle_info_nvx                                            = 1000030000
	image_view_address_properties_nvx                                     = 1000030001
	video_encode_h264_capabilities_khr                                    = 1000038000
	video_encode_h264_session_parameters_create_info_khr                  = 1000038001
	video_encode_h264_session_parameters_add_info_khr                     = 1000038002
	video_encode_h264_picture_info_khr                                    = 1000038003
	video_encode_h264_dpb_slot_info_khr                                   = 1000038004
	video_encode_h264_nalu_slice_info_khr                                 = 1000038005
	video_encode_h264_gop_remaining_frame_info_khr                        = 1000038006
	video_encode_h264_profile_info_khr                                    = 1000038007
	video_encode_h264_rate_control_info_khr                               = 1000038008
	video_encode_h264_rate_control_layer_info_khr                         = 1000038009
	video_encode_h264_session_create_info_khr                             = 1000038010
	video_encode_h264_quality_level_properties_khr                        = 1000038011
	video_encode_h264_session_parameters_get_info_khr                     = 1000038012
	video_encode_h264_session_parameters_feedback_info_khr                = 1000038013
	video_encode_h265_capabilities_khr                                    = 1000039000
	video_encode_h265_session_parameters_create_info_khr                  = 1000039001
	video_encode_h265_session_parameters_add_info_khr                     = 1000039002
	video_encode_h265_picture_info_khr                                    = 1000039003
	video_encode_h265_dpb_slot_info_khr                                   = 1000039004
	video_encode_h265_nalu_slice_segment_info_khr                         = 1000039005
	video_encode_h265_gop_remaining_frame_info_khr                        = 1000039006
	video_encode_h265_profile_info_khr                                    = 1000039007
	video_encode_h265_rate_control_info_khr                               = 1000039009
	video_encode_h265_rate_control_layer_info_khr                         = 1000039010
	video_encode_h265_session_create_info_khr                             = 1000039011
	video_encode_h265_quality_level_properties_khr                        = 1000039012
	video_encode_h265_session_parameters_get_info_khr                     = 1000039013
	video_encode_h265_session_parameters_feedback_info_khr                = 1000039014
	video_decode_h264_capabilities_khr                                    = 1000040000
	video_decode_h264_picture_info_khr                                    = 1000040001
	video_decode_h264_profile_info_khr                                    = 1000040003
	video_decode_h264_session_parameters_create_info_khr                  = 1000040004
	video_decode_h264_session_parameters_add_info_khr                     = 1000040005
	video_decode_h264_dpb_slot_info_khr                                   = 1000040006
	texture_lod_gather_format_properties_amd                              = 1000041000
	stream_descriptor_surface_create_info_ggp                             = 1000049000
	physical_device_corner_sampled_image_features_nv                      = 1000050000
	external_memory_image_create_info_nv                                  = 1000056000
	export_memory_allocate_info_nv                                        = 1000056001
	import_memory_win32_handle_info_nv                                    = 1000057000
	export_memory_win32_handle_info_nv                                    = 1000057001
	win32_keyed_mutex_acquire_release_info_nv                             = 1000058000
	validation_flags_ext                                                  = 1000061000
	vi_surface_create_info_nn                                             = 1000062000
	image_view_astc_decode_mode_ext                                       = 1000067000
	physical_device_astc_decode_features_ext                              = 1000067001
	import_memory_win32_handle_info_khr                                   = 1000073000
	export_memory_win32_handle_info_khr                                   = 1000073001
	memory_win32_handle_properties_khr                                    = 1000073002
	memory_get_win32_handle_info_khr                                      = 1000073003
	import_memory_fd_info_khr                                             = 1000074000
	memory_fd_properties_khr                                              = 1000074001
	memory_get_fd_info_khr                                                = 1000074002
	win32_keyed_mutex_acquire_release_info_khr                            = 1000075000
	import_semaphore_win32_handle_info_khr                                = 1000078000
	export_semaphore_win32_handle_info_khr                                = 1000078001
	d3d12_fence_submit_info_khr                                           = 1000078002
	semaphore_get_win32_handle_info_khr                                   = 1000078003
	import_semaphore_fd_info_khr                                          = 1000079000
	semaphore_get_fd_info_khr                                             = 1000079001
	command_buffer_inheritance_conditional_rendering_info_ext             = 1000081000
	physical_device_conditional_rendering_features_ext                    = 1000081001
	conditional_rendering_begin_info_ext                                  = 1000081002
	present_regions_khr                                                   = 1000084000
	pipeline_viewport_w_scaling_state_create_info_nv                      = 1000087000
	surface_capabilities2_ext                                             = 1000090000
	display_power_info_ext                                                = 1000091000
	device_event_info_ext                                                 = 1000091001
	display_event_info_ext                                                = 1000091002
	swapchain_counter_create_info_ext                                     = 1000091003
	present_times_info_google                                             = 1000092000
	physical_device_multiview_per_view_attributes_properties_nvx          = 1000097000
	multiview_per_view_attributes_info_nvx                                = 1000044009
	pipeline_viewport_swizzle_state_create_info_nv                        = 1000098000
	physical_device_discard_rectangle_properties_ext                      = 1000099000
	pipeline_discard_rectangle_state_create_info_ext                      = 1000099001
	physical_device_conservative_rasterization_properties_ext             = 1000101000
	pipeline_rasterization_conservative_state_create_info_ext             = 1000101001
	physical_device_depth_clip_enable_features_ext                        = 1000102000
	pipeline_rasterization_depth_clip_state_create_info_ext               = 1000102001
	hdr_metadata_ext                                                      = 1000105000
	physical_device_relaxed_line_rasterization_features_img               = 1000110000
	shared_present_surface_capabilities_khr                               = 1000111000
	import_fence_win32_handle_info_khr                                    = 1000114000
	export_fence_win32_handle_info_khr                                    = 1000114001
	fence_get_win32_handle_info_khr                                       = 1000114002
	import_fence_fd_info_khr                                              = 1000115000
	fence_get_fd_info_khr                                                 = 1000115001
	physical_device_performance_query_features_khr                        = 1000116000
	physical_device_performance_query_properties_khr                      = 1000116001
	query_pool_performance_create_info_khr                                = 1000116002
	performance_query_submit_info_khr                                     = 1000116003
	acquire_profiling_lock_info_khr                                       = 1000116004
	performance_counter_khr                                               = 1000116005
	performance_counter_description_khr                                   = 1000116006
	physical_device_surface_info2_khr                                     = 1000119000
	surface_capabilities2_khr                                             = 1000119001
	surface_format2_khr                                                   = 1000119002
	display_properties2_khr                                               = 1000121000
	display_plane_properties2_khr                                         = 1000121001
	display_mode_properties2_khr                                          = 1000121002
	display_plane_info2_khr                                               = 1000121003
	display_plane_capabilities2_khr                                       = 1000121004
	ios_surface_create_info_mvk                                           = 1000122000
	macos_surface_create_info_mvk                                         = 1000123000
	debug_utils_object_name_info_ext                                      = 1000128000
	debug_utils_object_tag_info_ext                                       = 1000128001
	debug_utils_label_ext                                                 = 1000128002
	debug_utils_messenger_callback_data_ext                               = 1000128003
	debug_utils_messenger_create_info_ext                                 = 1000128004
	android_hardware_buffer_usage_android                                 = 1000129000
	android_hardware_buffer_properties_android                            = 1000129001
	android_hardware_buffer_format_properties_android                     = 1000129002
	import_android_hardware_buffer_info_android                           = 1000129003
	memory_get_android_hardware_buffer_info_android                       = 1000129004
	external_format_android                                               = 1000129005
	android_hardware_buffer_format_properties2_android                    = 1000129006
	attachment_sample_count_info_amd                                      = 1000044008
	physical_device_shader_bfloat16_features_khr                          = 1000141000
	sample_locations_info_ext                                             = 1000143000
	render_pass_sample_locations_begin_info_ext                           = 1000143001
	pipeline_sample_locations_state_create_info_ext                       = 1000143002
	physical_device_sample_locations_properties_ext                       = 1000143003
	multisample_properties_ext                                            = 1000143004
	physical_device_blend_operation_advanced_features_ext                 = 1000148000
	physical_device_blend_operation_advanced_properties_ext               = 1000148001
	pipeline_color_blend_advanced_state_create_info_ext                   = 1000148002
	pipeline_coverage_to_color_state_create_info_nv                       = 1000149000
	write_descriptor_set_acceleration_structure_khr                       = 1000150007
	acceleration_structure_build_geometry_info_khr                        = 1000150000
	acceleration_structure_device_address_info_khr                        = 1000150002
	acceleration_structure_geometry_aabbs_data_khr                        = 1000150003
	acceleration_structure_geometry_instances_data_khr                    = 1000150004
	acceleration_structure_geometry_triangles_data_khr                    = 1000150005
	acceleration_structure_geometry_khr                                   = 1000150006
	acceleration_structure_version_info_khr                               = 1000150009
	copy_acceleration_structure_info_khr                                  = 1000150010
	copy_acceleration_structure_to_memory_info_khr                        = 1000150011
	copy_memory_to_acceleration_structure_info_khr                        = 1000150012
	physical_device_acceleration_structure_features_khr                   = 1000150013
	physical_device_acceleration_structure_properties_khr                 = 1000150014
	acceleration_structure_create_info_khr                                = 1000150017
	acceleration_structure_build_sizes_info_khr                           = 1000150020
	physical_device_ray_tracing_pipeline_features_khr                     = 1000347000
	physical_device_ray_tracing_pipeline_properties_khr                   = 1000347001
	ray_tracing_pipeline_create_info_khr                                  = 1000150015
	ray_tracing_shader_group_create_info_khr                              = 1000150016
	ray_tracing_pipeline_interface_create_info_khr                        = 1000150018
	physical_device_ray_query_features_khr                                = 1000348013
	pipeline_coverage_modulation_state_create_info_nv                     = 1000152000
	physical_device_shader_sm_builtins_features_nv                        = 1000154000
	physical_device_shader_sm_builtins_properties_nv                      = 1000154001
	drm_format_modifier_properties_list_ext                               = 1000158000
	physical_device_image_drm_format_modifier_info_ext                    = 1000158002
	image_drm_format_modifier_list_create_info_ext                        = 1000158003
	image_drm_format_modifier_explicit_create_info_ext                    = 1000158004
	image_drm_format_modifier_properties_ext                              = 1000158005
	drm_format_modifier_properties_list2_ext                              = 1000158006
	validation_cache_create_info_ext                                      = 1000160000
	shader_module_validation_cache_create_info_ext                        = 1000160001
	pipeline_viewport_shading_rate_image_state_create_info_nv             = 1000164000
	physical_device_shading_rate_image_features_nv                        = 1000164001
	physical_device_shading_rate_image_properties_nv                      = 1000164002
	pipeline_viewport_coarse_sample_order_state_create_info_nv            = 1000164005
	ray_tracing_pipeline_create_info_nv                                   = 1000165000
	acceleration_structure_create_info_nv                                 = 1000165001
	geometry_nv                                                           = 1000165003
	geometry_triangles_nv                                                 = 1000165004
	geometry_aabb_nv                                                      = 1000165005
	bind_acceleration_structure_memory_info_nv                            = 1000165006
	write_descriptor_set_acceleration_structure_nv                        = 1000165007
	acceleration_structure_memory_requirements_info_nv                    = 1000165008
	physical_device_ray_tracing_properties_nv                             = 1000165009
	ray_tracing_shader_group_create_info_nv                               = 1000165011
	acceleration_structure_info_nv                                        = 1000165012
	physical_device_representative_fragment_test_features_nv              = 1000166000
	pipeline_representative_fragment_test_state_create_info_nv            = 1000166001
	physical_device_image_view_image_format_info_ext                      = 1000170000
	filter_cubic_image_view_image_format_properties_ext                   = 1000170001
	import_memory_host_pointer_info_ext                                   = 1000178000
	memory_host_pointer_properties_ext                                    = 1000178001
	physical_device_external_memory_host_properties_ext                   = 1000178002
	physical_device_shader_clock_features_khr                             = 1000181000
	pipeline_compiler_control_create_info_amd                             = 1000183000
	physical_device_shader_core_properties_amd                            = 1000185000
	video_decode_h265_capabilities_khr                                    = 1000187000
	video_decode_h265_session_parameters_create_info_khr                  = 1000187001
	video_decode_h265_session_parameters_add_info_khr                     = 1000187002
	video_decode_h265_profile_info_khr                                    = 1000187003
	video_decode_h265_picture_info_khr                                    = 1000187004
	video_decode_h265_dpb_slot_info_khr                                   = 1000187005
	device_memory_overallocation_create_info_amd                          = 1000189000
	physical_device_vertex_attribute_divisor_properties_ext               = 1000190000
	present_frame_token_ggp                                               = 1000191000
	physical_device_mesh_shader_features_nv                               = 1000202000
	physical_device_mesh_shader_properties_nv                             = 1000202001
	physical_device_shader_image_footprint_features_nv                    = 1000204000
	pipeline_viewport_exclusive_scissor_state_create_info_nv              = 1000205000
	physical_device_exclusive_scissor_features_nv                         = 1000205002
	checkpoint_data_nv                                                    = 1000206000
	queue_family_checkpoint_properties_nv                                 = 1000206001
	queue_family_checkpoint_properties2_nv                                = 1000314008
	checkpoint_data2_nv                                                   = 1000314009
	physical_device_shader_integer_functions2_features_intel              = 1000209000
	query_pool_performance_query_create_info_intel                        = 1000210000
	initialize_performance_api_info_intel                                 = 1000210001
	performance_marker_info_intel                                         = 1000210002
	performance_stream_marker_info_intel                                  = 1000210003
	performance_override_info_intel                                       = 1000210004
	performance_configuration_acquire_info_intel                          = 1000210005
	physical_device_pci_bus_info_properties_ext                           = 1000212000
	display_native_hdr_surface_capabilities_amd                           = 1000213000
	swapchain_display_native_hdr_create_info_amd                          = 1000213001
	imagepipe_surface_create_info_fuchsia                                 = 1000214000
	metal_surface_create_info_ext                                         = 1000217000
	physical_device_fragment_density_map_features_ext                     = 1000218000
	physical_device_fragment_density_map_properties_ext                   = 1000218001
	render_pass_fragment_density_map_create_info_ext                      = 1000218002
	rendering_fragment_density_map_attachment_info_ext                    = 1000044007
	fragment_shading_rate_attachment_info_khr                             = 1000226000
	pipeline_fragment_shading_rate_state_create_info_khr                  = 1000226001
	physical_device_fragment_shading_rate_properties_khr                  = 1000226002
	physical_device_fragment_shading_rate_features_khr                    = 1000226003
	physical_device_fragment_shading_rate_khr                             = 1000226004
	rendering_fragment_shading_rate_attachment_info_khr                   = 1000044006
	physical_device_shader_core_properties2_amd                           = 1000227000
	physical_device_coherent_memory_features_amd                          = 1000229000
	physical_device_shader_image_atomic_int64_features_ext                = 1000234000
	physical_device_shader_quad_control_features_khr                      = 1000235000
	physical_device_memory_budget_properties_ext                          = 1000237000
	physical_device_memory_priority_features_ext                          = 1000238000
	memory_priority_allocate_info_ext                                     = 1000238001
	surface_protected_capabilities_khr                                    = 1000239000
	physical_device_dedicated_allocation_image_aliasing_features_nv       = 1000240000
	physical_device_buffer_device_address_features_ext                    = 1000244000
	buffer_device_address_create_info_ext                                 = 1000244002
	validation_features_ext                                               = 1000247000
	physical_device_present_wait_features_khr                             = 1000248000
	physical_device_cooperative_matrix_features_nv                        = 1000249000
	cooperative_matrix_properties_nv                                      = 1000249001
	physical_device_cooperative_matrix_properties_nv                      = 1000249002
	physical_device_coverage_reduction_mode_features_nv                   = 1000250000
	pipeline_coverage_reduction_state_create_info_nv                      = 1000250001
	framebuffer_mixed_samples_combination_nv                              = 1000250002
	physical_device_fragment_shader_interlock_features_ext                = 1000251000
	physical_device_ycbcr_image_arrays_features_ext                       = 1000252000
	physical_device_provoking_vertex_features_ext                         = 1000254000
	pipeline_rasterization_provoking_vertex_state_create_info_ext         = 1000254001
	physical_device_provoking_vertex_properties_ext                       = 1000254002
	surface_full_screen_exclusive_info_ext                                = 1000255000
	surface_capabilities_full_screen_exclusive_ext                        = 1000255002
	surface_full_screen_exclusive_win32_info_ext                          = 1000255001
	headless_surface_create_info_ext                                      = 1000256000
	physical_device_shader_atomic_float_features_ext                      = 1000260000
	physical_device_extended_dynamic_state_features_ext                   = 1000267000
	physical_device_pipeline_executable_properties_features_khr           = 1000269000
	pipeline_info_khr                                                     = 1000269001
	pipeline_executable_properties_khr                                    = 1000269002
	pipeline_executable_info_khr                                          = 1000269003
	pipeline_executable_statistic_khr                                     = 1000269004
	pipeline_executable_internal_representation_khr                       = 1000269005
	physical_device_map_memory_placed_features_ext                        = 1000272000
	physical_device_map_memory_placed_properties_ext                      = 1000272001
	memory_map_placed_info_ext                                            = 1000272002
	physical_device_shader_atomic_float2_features_ext                     = 1000273000
	physical_device_device_generated_commands_properties_nv               = 1000277000
	graphics_shader_group_create_info_nv                                  = 1000277001
	graphics_pipeline_shader_groups_create_info_nv                        = 1000277002
	indirect_commands_layout_token_nv                                     = 1000277003
	indirect_commands_layout_create_info_nv                               = 1000277004
	generated_commands_info_nv                                            = 1000277005
	generated_commands_memory_requirements_info_nv                        = 1000277006
	physical_device_device_generated_commands_features_nv                 = 1000277007
	physical_device_inherited_viewport_scissor_features_nv                = 1000278000
	command_buffer_inheritance_viewport_scissor_info_nv                   = 1000278001
	physical_device_texel_buffer_alignment_features_ext                   = 1000281000
	command_buffer_inheritance_render_pass_transform_info_qcom            = 1000282000
	render_pass_transform_begin_info_qcom                                 = 1000282001
	physical_device_depth_bias_control_features_ext                       = 1000283000
	depth_bias_info_ext                                                   = 1000283001
	depth_bias_representation_info_ext                                    = 1000283002
	physical_device_device_memory_report_features_ext                     = 1000284000
	device_device_memory_report_create_info_ext                           = 1000284001
	device_memory_report_callback_data_ext                                = 1000284002
	sampler_custom_border_color_create_info_ext                           = 1000287000
	physical_device_custom_border_color_properties_ext                    = 1000287001
	physical_device_custom_border_color_features_ext                      = 1000287002
	pipeline_library_create_info_khr                                      = 1000290000
	physical_device_present_barrier_features_nv                           = 1000292000
	surface_capabilities_present_barrier_nv                               = 1000292001
	swapchain_present_barrier_create_info_nv                              = 1000292002
	present_id_khr                                                        = 1000294000
	physical_device_present_id_features_khr                               = 1000294001
	video_encode_info_khr                                                 = 1000299000
	video_encode_rate_control_info_khr                                    = 1000299001
	video_encode_rate_control_layer_info_khr                              = 1000299002
	video_encode_capabilities_khr                                         = 1000299003
	video_encode_usage_info_khr                                           = 1000299004
	query_pool_video_encode_feedback_create_info_khr                      = 1000299005
	physical_device_video_encode_quality_level_info_khr                   = 1000299006
	video_encode_quality_level_properties_khr                             = 1000299007
	video_encode_quality_level_info_khr                                   = 1000299008
	video_encode_session_parameters_get_info_khr                          = 1000299009
	video_encode_session_parameters_feedback_info_khr                     = 1000299010
	physical_device_diagnostics_config_features_nv                        = 1000300000
	device_diagnostics_config_create_info_nv                              = 1000300001
	physical_device_tile_shading_features_qcom                            = 1000309000
	physical_device_tile_shading_properties_qcom                          = 1000309001
	render_pass_tile_shading_create_info_qcom                             = 1000309002
	per_tile_begin_info_qcom                                              = 1000309003
	per_tile_end_info_qcom                                                = 1000309004
	dispatch_tile_info_qcom                                               = 1000309005
	query_low_latency_support_nv                                          = 1000310000
	export_metal_object_create_info_ext                                   = 1000311000
	export_metal_objects_info_ext                                         = 1000311001
	export_metal_device_info_ext                                          = 1000311002
	export_metal_command_queue_info_ext                                   = 1000311003
	export_metal_buffer_info_ext                                          = 1000311004
	import_metal_buffer_info_ext                                          = 1000311005
	export_metal_texture_info_ext                                         = 1000311006
	import_metal_texture_info_ext                                         = 1000311007
	export_metal_io_surface_info_ext                                      = 1000311008
	import_metal_io_surface_info_ext                                      = 1000311009
	export_metal_shared_event_info_ext                                    = 1000311010
	import_metal_shared_event_info_ext                                    = 1000311011
	physical_device_descriptor_buffer_properties_ext                      = 1000316000
	physical_device_descriptor_buffer_density_map_properties_ext          = 1000316001
	physical_device_descriptor_buffer_features_ext                        = 1000316002
	descriptor_address_info_ext                                           = 1000316003
	descriptor_get_info_ext                                               = 1000316004
	buffer_capture_descriptor_data_info_ext                               = 1000316005
	image_capture_descriptor_data_info_ext                                = 1000316006
	image_view_capture_descriptor_data_info_ext                           = 1000316007
	sampler_capture_descriptor_data_info_ext                              = 1000316008
	opaque_capture_descriptor_data_create_info_ext                        = 1000316010
	descriptor_buffer_binding_info_ext                                    = 1000316011
	descriptor_buffer_binding_push_descriptor_buffer_handle_ext           = 1000316012
	acceleration_structure_capture_descriptor_data_info_ext               = 1000316009
	physical_device_graphics_pipeline_library_features_ext                = 1000320000
	physical_device_graphics_pipeline_library_properties_ext              = 1000320001
	graphics_pipeline_library_create_info_ext                             = 1000320002
	physical_device_shader_early_and_late_fragment_tests_features_amd     = 1000321000
	physical_device_fragment_shader_barycentric_features_khr              = 1000203000
	physical_device_fragment_shader_barycentric_properties_khr            = 1000322000
	physical_device_shader_subgroup_uniform_control_flow_features_khr     = 1000323000
	physical_device_fragment_shading_rate_enums_properties_nv             = 1000326000
	physical_device_fragment_shading_rate_enums_features_nv               = 1000326001
	pipeline_fragment_shading_rate_enum_state_create_info_nv              = 1000326002
	acceleration_structure_geometry_motion_triangles_data_nv              = 1000327000
	physical_device_ray_tracing_motion_blur_features_nv                   = 1000327001
	acceleration_structure_motion_info_nv                                 = 1000327002
	physical_device_mesh_shader_features_ext                              = 1000328000
	physical_device_mesh_shader_properties_ext                            = 1000328001
	physical_device_ycbcr2_plane444_formats_features_ext                  = 1000330000
	physical_device_fragment_density_map2_features_ext                    = 1000332000
	physical_device_fragment_density_map2_properties_ext                  = 1000332001
	copy_command_transform_info_qcom                                      = 1000333000
	physical_device_workgroup_memory_explicit_layout_features_khr         = 1000336000
	physical_device_image_compression_control_features_ext                = 1000338000
	image_compression_control_ext                                         = 1000338001
	image_compression_properties_ext                                      = 1000338004
	physical_device_attachment_feedback_loop_layout_features_ext          = 1000339000
	physical_device4444_formats_features_ext                              = 1000340000
	physical_device_fault_features_ext                                    = 1000341000
	device_fault_counts_ext                                               = 1000341001
	device_fault_info_ext                                                 = 1000341002
	physical_device_rgba10x6_formats_features_ext                         = 1000344000
	directfb_surface_create_info_ext                                      = 1000346000
	physical_device_vertex_input_dynamic_state_features_ext               = 1000352000
	vertex_input_binding_description2_ext                                 = 1000352001
	vertex_input_attribute_description2_ext                               = 1000352002
	physical_device_drm_properties_ext                                    = 1000353000
	physical_device_address_binding_report_features_ext                   = 1000354000
	device_address_binding_callback_data_ext                              = 1000354001
	physical_device_depth_clip_control_features_ext                       = 1000355000
	pipeline_viewport_depth_clip_control_create_info_ext                  = 1000355001
	physical_device_primitive_topology_list_restart_features_ext          = 1000356000
	import_memory_zircon_handle_info_fuchsia                              = 1000364000
	memory_zircon_handle_properties_fuchsia                               = 1000364001
	memory_get_zircon_handle_info_fuchsia                                 = 1000364002
	import_semaphore_zircon_handle_info_fuchsia                           = 1000365000
	semaphore_get_zircon_handle_info_fuchsia                              = 1000365001
	buffer_collection_create_info_fuchsia                                 = 1000366000
	import_memory_buffer_collection_fuchsia                               = 1000366001
	buffer_collection_image_create_info_fuchsia                           = 1000366002
	buffer_collection_properties_fuchsia                                  = 1000366003
	buffer_constraints_info_fuchsia                                       = 1000366004
	buffer_collection_buffer_create_info_fuchsia                          = 1000366005
	image_constraints_info_fuchsia                                        = 1000366006
	image_format_constraints_info_fuchsia                                 = 1000366007
	sysmem_color_space_fuchsia                                            = 1000366008
	buffer_collection_constraints_info_fuchsia                            = 1000366009
	subpass_shading_pipeline_create_info_huawei                           = 1000369000
	physical_device_subpass_shading_features_huawei                       = 1000369001
	physical_device_subpass_shading_properties_huawei                     = 1000369002
	physical_device_invocation_mask_features_huawei                       = 1000370000
	memory_get_remote_address_info_nv                                     = 1000371000
	physical_device_external_memory_rdma_features_nv                      = 1000371001
	pipeline_properties_identifier_ext                                    = 1000372000
	physical_device_pipeline_properties_features_ext                      = 1000372001
	physical_device_frame_boundary_features_ext                           = 1000375000
	frame_boundary_ext                                                    = 1000375001
	physical_device_multisampled_render_to_single_sampled_features_ext    = 1000376000
	subpass_resolve_performance_query_ext                                 = 1000376001
	multisampled_render_to_single_sampled_info_ext                        = 1000376002
	physical_device_extended_dynamic_state2_features_ext                  = 1000377000
	screen_surface_create_info_qnx                                        = 1000378000
	physical_device_color_write_enable_features_ext                       = 1000381000
	pipeline_color_write_create_info_ext                                  = 1000381001
	physical_device_primitives_generated_query_features_ext               = 1000382000
	physical_device_ray_tracing_maintenance1_features_khr                 = 1000386000
	physical_device_shader_untyped_pointers_features_khr                  = 1000387000
	physical_device_video_encode_rgb_conversion_features_valve            = 1000390000
	video_encode_rgb_conversion_capabilities_valve                        = 1000390001
	video_encode_profile_rgb_conversion_info_valve                        = 1000390002
	video_encode_session_rgb_conversion_create_info_valve                 = 1000390003
	physical_device_image_view_min_lod_features_ext                       = 1000391000
	image_view_min_lod_create_info_ext                                    = 1000391001
	physical_device_multi_draw_features_ext                               = 1000392000
	physical_device_multi_draw_properties_ext                             = 1000392001
	physical_device_image2d_view_of3d_features_ext                        = 1000393000
	physical_device_shader_tile_image_features_ext                        = 1000395000
	physical_device_shader_tile_image_properties_ext                      = 1000395001
	micromap_build_info_ext                                               = 1000396000
	micromap_version_info_ext                                             = 1000396001
	copy_micromap_info_ext                                                = 1000396002
	copy_micromap_to_memory_info_ext                                      = 1000396003
	copy_memory_to_micromap_info_ext                                      = 1000396004
	physical_device_opacity_micromap_features_ext                         = 1000396005
	physical_device_opacity_micromap_properties_ext                       = 1000396006
	micromap_create_info_ext                                              = 1000396007
	micromap_build_sizes_info_ext                                         = 1000396008
	acceleration_structure_triangles_opacity_micromap_ext                 = 1000396009
	physical_device_cluster_culling_shader_features_huawei                = 1000404000
	physical_device_cluster_culling_shader_properties_huawei              = 1000404001
	physical_device_cluster_culling_shader_vrs_features_huawei            = 1000404002
	physical_device_border_color_swizzle_features_ext                     = 1000411000
	sampler_border_color_component_mapping_create_info_ext                = 1000411001
	physical_device_pageable_device_local_memory_features_ext             = 1000412000
	physical_device_shader_core_properties_arm                            = 1000415000
	device_queue_shader_core_control_create_info_arm                      = 1000417000
	physical_device_scheduling_controls_features_arm                      = 1000417001
	physical_device_scheduling_controls_properties_arm                    = 1000417002
	physical_device_image_sliced_view_of3d_features_ext                   = 1000418000
	image_view_sliced_create_info_ext                                     = 1000418001
	physical_device_descriptor_set_host_mapping_features_valve            = 1000420000
	descriptor_set_binding_reference_valve                                = 1000420001
	descriptor_set_layout_host_mapping_info_valve                         = 1000420002
	physical_device_non_seamless_cube_map_features_ext                    = 1000422000
	physical_device_render_pass_striped_features_arm                      = 1000424000
	physical_device_render_pass_striped_properties_arm                    = 1000424001
	render_pass_stripe_begin_info_arm                                     = 1000424002
	render_pass_stripe_info_arm                                           = 1000424003
	render_pass_stripe_submit_info_arm                                    = 1000424004
	physical_device_copy_memory_indirect_features_nv                      = 1000426000
	physical_device_device_generated_commands_compute_features_nv         = 1000428000
	compute_pipeline_indirect_buffer_info_nv                              = 1000428001
	pipeline_indirect_device_address_info_nv                              = 1000428002
	physical_device_ray_tracing_linear_swept_spheres_features_nv          = 1000429008
	acceleration_structure_geometry_linear_swept_spheres_data_nv          = 1000429009
	acceleration_structure_geometry_spheres_data_nv                       = 1000429010
	physical_device_linear_color_attachment_features_nv                   = 1000430000
	physical_device_shader_maximal_reconvergence_features_khr             = 1000434000
	physical_device_image_compression_control_swapchain_features_ext      = 1000437000
	physical_device_image_processing_features_qcom                        = 1000440000
	physical_device_image_processing_properties_qcom                      = 1000440001
	image_view_sample_weight_create_info_qcom                             = 1000440002
	physical_device_nested_command_buffer_features_ext                    = 1000451000
	physical_device_nested_command_buffer_properties_ext                  = 1000451001
	external_memory_acquire_unmodified_ext                                = 1000453000
	physical_device_extended_dynamic_state3_features_ext                  = 1000455000
	physical_device_extended_dynamic_state3_properties_ext                = 1000455001
	physical_device_subpass_merge_feedback_features_ext                   = 1000458000
	render_pass_creation_control_ext                                      = 1000458001
	render_pass_creation_feedback_create_info_ext                         = 1000458002
	render_pass_subpass_feedback_create_info_ext                          = 1000458003
	direct_driver_loading_info_lunarg                                     = 1000459000
	direct_driver_loading_list_lunarg                                     = 1000459001
	tensor_create_info_arm                                                = 1000460000
	tensor_view_create_info_arm                                           = 1000460001
	bind_tensor_memory_info_arm                                           = 1000460002
	write_descriptor_set_tensor_arm                                       = 1000460003
	physical_device_tensor_properties_arm                                 = 1000460004
	tensor_format_properties_arm                                          = 1000460005
	tensor_description_arm                                                = 1000460006
	tensor_memory_requirements_info_arm                                   = 1000460007
	tensor_memory_barrier_arm                                             = 1000460008
	physical_device_tensor_features_arm                                   = 1000460009
	device_tensor_memory_requirements_arm                                 = 1000460010
	copy_tensor_info_arm                                                  = 1000460011
	tensor_copy_arm                                                       = 1000460012
	tensor_dependency_info_arm                                            = 1000460013
	memory_dedicated_allocate_info_tensor_arm                             = 1000460014
	physical_device_external_tensor_info_arm                              = 1000460015
	external_tensor_properties_arm                                        = 1000460016
	external_memory_tensor_create_info_arm                                = 1000460017
	physical_device_descriptor_buffer_tensor_features_arm                 = 1000460018
	physical_device_descriptor_buffer_tensor_properties_arm               = 1000460019
	descriptor_get_tensor_info_arm                                        = 1000460020
	tensor_capture_descriptor_data_info_arm                               = 1000460021
	tensor_view_capture_descriptor_data_info_arm                          = 1000460022
	frame_boundary_tensors_arm                                            = 1000460023
	physical_device_shader_module_identifier_features_ext                 = 1000462000
	physical_device_shader_module_identifier_properties_ext               = 1000462001
	pipeline_shader_stage_module_identifier_create_info_ext               = 1000462002
	shader_module_identifier_ext                                          = 1000462003
	physical_device_rasterization_order_attachment_access_features_ext    = 1000342000
	physical_device_optical_flow_features_nv                              = 1000464000
	physical_device_optical_flow_properties_nv                            = 1000464001
	optical_flow_image_format_info_nv                                     = 1000464002
	optical_flow_image_format_properties_nv                               = 1000464003
	optical_flow_session_create_info_nv                                   = 1000464004
	optical_flow_execute_info_nv                                          = 1000464005
	optical_flow_session_create_private_data_info_nv                      = 1000464010
	physical_device_legacy_dithering_features_ext                         = 1000465000
	physical_device_external_format_resolve_features_android              = 1000468000
	physical_device_external_format_resolve_properties_android            = 1000468001
	android_hardware_buffer_format_resolve_properties_android             = 1000468002
	physical_device_anti_lag_features_amd                                 = 1000476000
	anti_lag_data_amd                                                     = 1000476001
	anti_lag_presentation_info_amd                                        = 1000476002
	surface_capabilities_present_id2_khr                                  = 1000479000
	present_id2_khr                                                       = 1000479001
	physical_device_present_id2_features_khr                              = 1000479002
	surface_capabilities_present_wait2_khr                                = 1000480000
	physical_device_present_wait2_features_khr                            = 1000480001
	present_wait2_info_khr                                                = 1000480002
	physical_device_ray_tracing_position_fetch_features_khr               = 1000481000
	physical_device_shader_object_features_ext                            = 1000482000
	physical_device_shader_object_properties_ext                          = 1000482001
	shader_create_info_ext                                                = 1000482002
	physical_device_pipeline_binary_features_khr                          = 1000483000
	pipeline_binary_create_info_khr                                       = 1000483001
	pipeline_binary_info_khr                                              = 1000483002
	pipeline_binary_key_khr                                               = 1000483003
	physical_device_pipeline_binary_properties_khr                        = 1000483004
	release_captured_pipeline_data_info_khr                               = 1000483005
	pipeline_binary_data_info_khr                                         = 1000483006
	pipeline_create_info_khr                                              = 1000483007
	device_pipeline_binary_internal_cache_control_khr                     = 1000483008
	pipeline_binary_handles_info_khr                                      = 1000483009
	physical_device_tile_properties_features_qcom                         = 1000484000
	tile_properties_qcom                                                  = 1000484001
	physical_device_amigo_profiling_features_sec                          = 1000485000
	amigo_profiling_submit_info_sec                                       = 1000485001
	surface_present_mode_khr                                              = 1000274000
	surface_present_scaling_capabilities_khr                              = 1000274001
	surface_present_mode_compatibility_khr                                = 1000274002
	physical_device_swapchain_maintenance1_features_khr                   = 1000275000
	swapchain_present_fence_info_khr                                      = 1000275001
	swapchain_present_modes_create_info_khr                               = 1000275002
	swapchain_present_mode_info_khr                                       = 1000275003
	swapchain_present_scaling_create_info_khr                             = 1000275004
	release_swapchain_images_info_khr                                     = 1000275005
	physical_device_multiview_per_view_viewports_features_qcom            = 1000488000
	physical_device_ray_tracing_invocation_reorder_features_nv            = 1000490000
	physical_device_ray_tracing_invocation_reorder_properties_nv          = 1000490001
	physical_device_cooperative_vector_features_nv                        = 1000491000
	physical_device_cooperative_vector_properties_nv                      = 1000491001
	cooperative_vector_properties_nv                                      = 1000491002
	convert_cooperative_vector_matrix_info_nv                             = 1000491004
	physical_device_extended_sparse_address_space_features_nv             = 1000492000
	physical_device_extended_sparse_address_space_properties_nv           = 1000492001
	physical_device_mutable_descriptor_type_features_ext                  = 1000351000
	mutable_descriptor_type_create_info_ext                               = 1000351002
	physical_device_legacy_vertex_attributes_features_ext                 = 1000495000
	physical_device_legacy_vertex_attributes_properties_ext               = 1000495001
	layer_settings_create_info_ext                                        = 1000496000
	physical_device_shader_core_builtins_features_arm                     = 1000497000
	physical_device_shader_core_builtins_properties_arm                   = 1000497001
	physical_device_pipeline_library_group_handles_features_ext           = 1000498000
	physical_device_dynamic_rendering_unused_attachments_features_ext     = 1000499000
	latency_sleep_mode_info_nv                                            = 1000505000
	latency_sleep_info_nv                                                 = 1000505001
	set_latency_marker_info_nv                                            = 1000505002
	get_latency_marker_info_nv                                            = 1000505003
	latency_timings_frame_report_nv                                       = 1000505004
	latency_submission_present_id_nv                                      = 1000505005
	out_of_band_queue_type_info_nv                                        = 1000505006
	swapchain_latency_create_info_nv                                      = 1000505007
	latency_surface_capabilities_nv                                       = 1000505008
	physical_device_cooperative_matrix_features_khr                       = 1000506000
	cooperative_matrix_properties_khr                                     = 1000506001
	physical_device_cooperative_matrix_properties_khr                     = 1000506002
	data_graph_pipeline_create_info_arm                                   = 1000507000
	data_graph_pipeline_session_create_info_arm                           = 1000507001
	data_graph_pipeline_resource_info_arm                                 = 1000507002
	data_graph_pipeline_constant_arm                                      = 1000507003
	data_graph_pipeline_session_memory_requirements_info_arm              = 1000507004
	bind_data_graph_pipeline_session_memory_info_arm                      = 1000507005
	physical_device_data_graph_features_arm                               = 1000507006
	data_graph_pipeline_shader_module_create_info_arm                     = 1000507007
	data_graph_pipeline_property_query_result_arm                         = 1000507008
	data_graph_pipeline_info_arm                                          = 1000507009
	data_graph_pipeline_compiler_control_create_info_arm                  = 1000507010
	data_graph_pipeline_session_bind_point_requirements_info_arm          = 1000507011
	data_graph_pipeline_session_bind_point_requirement_arm                = 1000507012
	data_graph_pipeline_identifier_create_info_arm                        = 1000507013
	data_graph_pipeline_dispatch_info_arm                                 = 1000507014
	data_graph_processing_engine_create_info_arm                          = 1000507016
	queue_family_data_graph_processing_engine_properties_arm              = 1000507017
	queue_family_data_graph_properties_arm                                = 1000507018
	physical_device_queue_family_data_graph_processing_engine_info_arm    = 1000507019
	data_graph_pipeline_constant_tensor_semi_structured_sparsity_info_arm = 1000507015
	physical_device_multiview_per_view_render_areas_features_qcom         = 1000510000
	multiview_per_view_render_areas_render_pass_begin_info_qcom           = 1000510001
	physical_device_compute_shader_derivatives_features_khr               = 1000201000
	physical_device_compute_shader_derivatives_properties_khr             = 1000511000
	video_decode_av1_capabilities_khr                                     = 1000512000
	video_decode_av1_picture_info_khr                                     = 1000512001
	video_decode_av1_profile_info_khr                                     = 1000512003
	video_decode_av1_session_parameters_create_info_khr                   = 1000512004
	video_decode_av1_dpb_slot_info_khr                                    = 1000512005
	video_encode_av1_capabilities_khr                                     = 1000513000
	video_encode_av1_session_parameters_create_info_khr                   = 1000513001
	video_encode_av1_picture_info_khr                                     = 1000513002
	video_encode_av1_dpb_slot_info_khr                                    = 1000513003
	physical_device_video_encode_av1_features_khr                         = 1000513004
	video_encode_av1_profile_info_khr                                     = 1000513005
	video_encode_av1_rate_control_info_khr                                = 1000513006
	video_encode_av1_rate_control_layer_info_khr                          = 1000513007
	video_encode_av1_quality_level_properties_khr                         = 1000513008
	video_encode_av1_session_create_info_khr                              = 1000513009
	video_encode_av1_gop_remaining_frame_info_khr                         = 1000513010
	physical_device_video_decode_vp9_features_khr                         = 1000514000
	video_decode_vp9_capabilities_khr                                     = 1000514001
	video_decode_vp9_picture_info_khr                                     = 1000514002
	video_decode_vp9_profile_info_khr                                     = 1000514003
	physical_device_video_maintenance1_features_khr                       = 1000515000
	video_inline_query_info_khr                                           = 1000515001
	physical_device_per_stage_descriptor_set_features_nv                  = 1000516000
	physical_device_image_processing2_features_qcom                       = 1000518000
	physical_device_image_processing2_properties_qcom                     = 1000518001
	sampler_block_match_window_create_info_qcom                           = 1000518002
	sampler_cubic_weights_create_info_qcom                                = 1000519000
	physical_device_cubic_weights_features_qcom                           = 1000519001
	blit_image_cubic_weights_info_qcom                                    = 1000519002
	physical_device_ycbcr_degamma_features_qcom                           = 1000520000
	sampler_ycbcr_conversion_ycbcr_degamma_create_info_qcom               = 1000520001
	physical_device_cubic_clamp_features_qcom                             = 1000521000
	physical_device_attachment_feedback_loop_dynamic_state_features_ext   = 1000524000
	physical_device_unified_image_layouts_features_khr                    = 1000527000
	attachment_feedback_loop_info_ext                                     = 1000527001
	screen_buffer_properties_qnx                                          = 1000529000
	screen_buffer_format_properties_qnx                                   = 1000529001
	import_screen_buffer_info_qnx                                         = 1000529002
	external_format_qnx                                                   = 1000529003
	physical_device_external_memory_screen_buffer_features_qnx            = 1000529004
	physical_device_layered_driver_properties_msft                        = 1000530000
	calibrated_timestamp_info_khr                                         = 1000184000
	set_descriptor_buffer_offsets_info_ext                                = 1000545007
	bind_descriptor_buffer_embedded_samplers_info_ext                     = 1000545008
	physical_device_descriptor_pool_overallocation_features_nv            = 1000546000
	physical_device_tile_memory_heap_features_qcom                        = 1000547000
	physical_device_tile_memory_heap_properties_qcom                      = 1000547001
	tile_memory_requirements_qcom                                         = 1000547002
	tile_memory_bind_info_qcom                                            = 1000547003
	tile_memory_size_info_qcom                                            = 1000547004
	physical_device_copy_memory_indirect_features_khr                     = 1000549000
	physical_device_copy_memory_indirect_properties_khr                   = 1000426001
	copy_memory_indirect_info_khr                                         = 1000549002
	copy_memory_to_image_indirect_info_khr                                = 1000549003
	physical_device_memory_decompression_features_ext                     = 1000427000
	physical_device_memory_decompression_properties_ext                   = 1000427001
	decompress_memory_info_ext                                            = 1000550002
	display_surface_stereo_create_info_nv                                 = 1000551000
	display_mode_stereo_properties_nv                                     = 1000551001
	video_encode_intra_refresh_capabilities_khr                           = 1000552000
	video_encode_session_intra_refresh_create_info_khr                    = 1000552001
	video_encode_intra_refresh_info_khr                                   = 1000552002
	video_reference_intra_refresh_info_khr                                = 1000552003
	physical_device_video_encode_intra_refresh_features_khr               = 1000552004
	video_encode_quantization_map_capabilities_khr                        = 1000553000
	video_format_quantization_map_properties_khr                          = 1000553001
	video_encode_quantization_map_info_khr                                = 1000553002
	video_encode_quantization_map_session_parameters_create_info_khr      = 1000553005
	physical_device_video_encode_quantization_map_features_khr            = 1000553009
	video_encode_h264_quantization_map_capabilities_khr                   = 1000553003
	video_encode_h265_quantization_map_capabilities_khr                   = 1000553004
	video_format_h265_quantization_map_properties_khr                     = 1000553006
	video_encode_av1_quantization_map_capabilities_khr                    = 1000553007
	video_format_av1_quantization_map_properties_khr                      = 1000553008
	physical_device_raw_access_chains_features_nv                         = 1000555000
	external_compute_queue_device_create_info_nv                          = 1000556000
	external_compute_queue_create_info_nv                                 = 1000556001
	external_compute_queue_data_params_nv                                 = 1000556002
	physical_device_external_compute_queue_properties_nv                  = 1000556003
	physical_device_shader_relaxed_extended_instruction_features_khr      = 1000558000
	physical_device_command_buffer_inheritance_features_nv                = 1000559000
	physical_device_maintenance7_features_khr                             = 1000562000
	physical_device_maintenance7_properties_khr                           = 1000562001
	physical_device_layered_api_properties_list_khr                       = 1000562002
	physical_device_layered_api_properties_khr                            = 1000562003
	physical_device_layered_api_vulkan_properties_khr                     = 1000562004
	physical_device_shader_atomic_float16_vector_features_nv              = 1000563000
	physical_device_shader_replicated_composites_features_ext             = 1000564000
	physical_device_shader_float8_features_ext                            = 1000567000
	physical_device_ray_tracing_validation_features_nv                    = 1000568000
	physical_device_cluster_acceleration_structure_features_nv            = 1000569000
	physical_device_cluster_acceleration_structure_properties_nv          = 1000569001
	cluster_acceleration_structure_clusters_bottom_level_input_nv         = 1000569002
	cluster_acceleration_structure_triangle_cluster_input_nv              = 1000569003
	cluster_acceleration_structure_move_objects_input_nv                  = 1000569004
	cluster_acceleration_structure_input_info_nv                          = 1000569005
	cluster_acceleration_structure_commands_info_nv                       = 1000569006
	ray_tracing_pipeline_cluster_acceleration_structure_create_info_nv    = 1000569007
	physical_device_partitioned_acceleration_structure_features_nv        = 1000570000
	physical_device_partitioned_acceleration_structure_properties_nv      = 1000570001
	write_descriptor_set_partitioned_acceleration_structure_nv            = 1000570002
	partitioned_acceleration_structure_instances_input_nv                 = 1000570003
	build_partitioned_acceleration_structure_info_nv                      = 1000570004
	partitioned_acceleration_structure_flags_nv                           = 1000570005
	physical_device_device_generated_commands_features_ext                = 1000572000
	physical_device_device_generated_commands_properties_ext              = 1000572001
	generated_commands_memory_requirements_info_ext                       = 1000572002
	indirect_execution_set_create_info_ext                                = 1000572003
	generated_commands_info_ext                                           = 1000572004
	indirect_commands_layout_create_info_ext                              = 1000572006
	indirect_commands_layout_token_ext                                    = 1000572007
	write_indirect_execution_set_pipeline_ext                             = 1000572008
	write_indirect_execution_set_shader_ext                               = 1000572009
	indirect_execution_set_pipeline_info_ext                              = 1000572010
	indirect_execution_set_shader_info_ext                                = 1000572011
	indirect_execution_set_shader_layout_info_ext                         = 1000572012
	generated_commands_pipeline_info_ext                                  = 1000572013
	generated_commands_shader_info_ext                                    = 1000572014
	physical_device_maintenance8_features_khr                             = 1000574000
	memory_barrier_access_flags3_khr                                      = 1000574002
	physical_device_image_alignment_control_features_mesa                 = 1000575000
	physical_device_image_alignment_control_properties_mesa               = 1000575001
	image_alignment_control_create_info_mesa                              = 1000575002
	physical_device_shader_fma_features_khr                               = 1000579000
	physical_device_depth_clamp_control_features_ext                      = 1000582000
	pipeline_viewport_depth_clamp_control_create_info_ext                 = 1000582001
	physical_device_maintenance9_features_khr                             = 1000584000
	physical_device_maintenance9_properties_khr                           = 1000584001
	queue_family_ownership_transfer_properties_khr                        = 1000584002
	physical_device_video_maintenance2_features_khr                       = 1000586000
	video_decode_h264_inline_session_parameters_info_khr                  = 1000586001
	video_decode_h265_inline_session_parameters_info_khr                  = 1000586002
	video_decode_av1_inline_session_parameters_info_khr                   = 1000586003
	surface_create_info_ohos                                              = 1000685000
	native_buffer_ohos                                                    = 1000453001
	swapchain_image_create_info_ohos                                      = 1000453002
	physical_device_presentation_properties_ohos                          = 1000453003
	physical_device_hdr_vivid_features_huawei                             = 1000590000
	hdr_vivid_dynamic_metadata_huawei                                     = 1000590001
	physical_device_cooperative_matrix2_features_nv                       = 1000593000
	cooperative_matrix_flexible_dimensions_properties_nv                  = 1000593001
	physical_device_cooperative_matrix2_properties_nv                     = 1000593002
	physical_device_pipeline_opacity_micromap_features_arm                = 1000596000
	import_memory_metal_handle_info_ext                                   = 1000602000
	memory_metal_handle_properties_ext                                    = 1000602001
	memory_get_metal_handle_info_ext                                      = 1000602002
	physical_device_depth_clamp_zero_one_features_khr                     = 1000421000
	physical_device_vertex_attribute_robustness_features_ext              = 1000608000
	physical_device_format_pack_features_arm                              = 1000609000
	physical_device_fragment_density_map_layered_features_valve           = 1000611000
	physical_device_fragment_density_map_layered_properties_valve         = 1000611001
	pipeline_fragment_density_map_layered_create_info_valve               = 1000611002
	physical_device_robustness2_features_khr                              = 1000286000
	physical_device_robustness2_properties_khr                            = 1000286001
	physical_device_fragment_density_map_offset_features_ext              = 1000425000
	physical_device_fragment_density_map_offset_properties_ext            = 1000425001
	render_pass_fragment_density_map_offset_end_info_ext                  = 1000425002
	physical_device_zero_initialize_device_memory_features_ext            = 1000620000
	physical_device_present_mode_fifo_latest_ready_features_khr           = 1000361000
	physical_device_shader64_bit_indexing_features_ext                    = 1000627000
	physical_device_maintenance10_features_khr                            = 1000630000
	physical_device_maintenance10_properties_khr                          = 1000630001
	rendering_attachment_flags_info_khr                                   = 1000630002
	rendering_end_info_khr                                                = 1000619003
	resolve_image_mode_info_khr                                           = 1000630004
	physical_device_pipeline_cache_incremental_mode_features_sec          = 1000637000
	physical_device_shader_uniform_buffer_unsized_array_features_ext      = 1000642000
	max_enum                                                              = max_int
}

pub enum ImageLayout as u32 {
	undefined                                    = 0
	general                                      = 1
	color_attachment_optimal                     = 2
	depth_stencil_attachment_optimal             = 3
	depth_stencil_read_only_optimal              = 4
	shader_read_only_optimal                     = 5
	transfer_src_optimal                         = 6
	transfer_dst_optimal                         = 7
	preinitialized                               = 8
	depth_read_only_stencil_attachment_optimal   = 1000117000
	depth_attachment_stencil_read_only_optimal   = 1000117001
	depth_attachment_optimal                     = 1000241000
	depth_read_only_optimal                      = 1000241001
	stencil_attachment_optimal                   = 1000241002
	stencil_read_only_optimal                    = 1000241003
	read_only_optimal                            = 1000314000
	attachment_optimal                           = 1000314001
	rendering_local_read                         = 1000232000
	present_src_khr                              = 1000001002
	video_decode_dst_khr                         = 1000024000
	video_decode_src_khr                         = 1000024001
	video_decode_dpb_khr                         = 1000024002
	shared_present_khr                           = 1000111000
	fragment_density_map_optimal_ext             = 1000218000
	fragment_shading_rate_attachment_optimal_khr = 1000164003
	video_encode_dst_khr                         = 1000299000
	video_encode_src_khr                         = 1000299001
	video_encode_dpb_khr                         = 1000299002
	attachment_feedback_loop_optimal_ext         = 1000339000
	tensor_aliasing_arm                          = 1000460000
	video_encode_quantization_map_khr            = 1000553000
	zero_initialized_ext                         = 1000620000
	max_enum                                     = max_int
}

pub enum ObjectType as u32 {
	unknown                         = 0
	instance                        = 1
	physical_device                 = 2
	device                          = 3
	queue                           = 4
	semaphore                       = 5
	command_buffer                  = 6
	fence                           = 7
	device_memory                   = 8
	buffer                          = 9
	image                           = 10
	event                           = 11
	query_pool                      = 12
	buffer_view                     = 13
	image_view                      = 14
	shader_module                   = 15
	pipeline_cache                  = 16
	pipeline_layout                 = 17
	render_pass                     = 18
	pipeline                        = 19
	descriptor_set_layout           = 20
	sampler                         = 21
	descriptor_pool                 = 22
	descriptor_set                  = 23
	framebuffer                     = 24
	command_pool                    = 25
	descriptor_update_template      = 1000085000
	sampler_ycbcr_conversion        = 1000156000
	private_data_slot               = 1000295000
	surface_khr                     = 1000000000
	swapchain_khr                   = 1000001000
	display_khr                     = 1000002000
	display_mode_khr                = 1000002001
	debug_report_callback_ext       = 1000011000
	video_session_khr               = 1000023000
	video_session_parameters_khr    = 1000023001
	cu_module_nvx                   = 1000029000
	cu_function_nvx                 = 1000029001
	debug_utils_messenger_ext       = 1000128000
	acceleration_structure_khr      = 1000150000
	validation_cache_ext            = 1000160000
	acceleration_structure_nv       = 1000165000
	performance_configuration_intel = 1000210000
	deferred_operation_khr          = 1000268000
	indirect_commands_layout_nv     = 1000277000
	buffer_collection_fuchsia       = 1000366000
	micromap_ext                    = 1000396000
	tensor_arm                      = 1000460000
	tensor_view_arm                 = 1000460001
	optical_flow_session_nv         = 1000464000
	shader_ext                      = 1000482000
	pipeline_binary_khr             = 1000483000
	data_graph_pipeline_session_arm = 1000507000
	external_compute_queue_nv       = 1000556000
	indirect_commands_layout_ext    = 1000572000
	indirect_execution_set_ext      = 1000572001
	max_enum                        = max_int
}

pub enum VendorId as u32 {
	khronos  = u32(0x10000)
	viv      = u32(0x10001)
	vsi      = u32(0x10002)
	kazan    = u32(0x10003)
	codeplay = u32(0x10004)
	mesa     = u32(0x10005)
	pocl     = u32(0x10006)
	mobileye = u32(0x10007)
	max_enum = max_int
}

pub enum SystemAllocationScope as u32 {
	command  = 0
	object   = 1
	cache    = 2
	device   = 3
	instance = 4
	max_enum = max_int
}

pub enum InternalAllocationType as u32 {
	executable = 0
	max_enum   = max_int
}

pub enum Format as u32 {
	undefined                                   = 0
	r4g4_unorm_pack8                            = 1
	r4g4b4a4_unorm_pack16                       = 2
	b4g4r4a4_unorm_pack16                       = 3
	r5g6b5_unorm_pack16                         = 4
	b5g6r5_unorm_pack16                         = 5
	r5g5b5a1_unorm_pack16                       = 6
	b5g5r5a1_unorm_pack16                       = 7
	a1r5g5b5_unorm_pack16                       = 8
	r8_unorm                                    = 9
	r8_snorm                                    = 10
	r8_uscaled                                  = 11
	r8_sscaled                                  = 12
	r8_uint                                     = 13
	r8_sint                                     = 14
	r8_srgb                                     = 15
	r8g8_unorm                                  = 16
	r8g8_snorm                                  = 17
	r8g8_uscaled                                = 18
	r8g8_sscaled                                = 19
	r8g8_uint                                   = 20
	r8g8_sint                                   = 21
	r8g8_srgb                                   = 22
	r8g8b8_unorm                                = 23
	r8g8b8_snorm                                = 24
	r8g8b8_uscaled                              = 25
	r8g8b8_sscaled                              = 26
	r8g8b8_uint                                 = 27
	r8g8b8_sint                                 = 28
	r8g8b8_srgb                                 = 29
	b8g8r8_unorm                                = 30
	b8g8r8_snorm                                = 31
	b8g8r8_uscaled                              = 32
	b8g8r8_sscaled                              = 33
	b8g8r8_uint                                 = 34
	b8g8r8_sint                                 = 35
	b8g8r8_srgb                                 = 36
	r8g8b8a8_unorm                              = 37
	r8g8b8a8_snorm                              = 38
	r8g8b8a8_uscaled                            = 39
	r8g8b8a8_sscaled                            = 40
	r8g8b8a8_uint                               = 41
	r8g8b8a8_sint                               = 42
	r8g8b8a8_srgb                               = 43
	b8g8r8a8_unorm                              = 44
	b8g8r8a8_snorm                              = 45
	b8g8r8a8_uscaled                            = 46
	b8g8r8a8_sscaled                            = 47
	b8g8r8a8_uint                               = 48
	b8g8r8a8_sint                               = 49
	b8g8r8a8_srgb                               = 50
	a8b8g8r8_unorm_pack32                       = 51
	a8b8g8r8_snorm_pack32                       = 52
	a8b8g8r8_uscaled_pack32                     = 53
	a8b8g8r8_sscaled_pack32                     = 54
	a8b8g8r8_uint_pack32                        = 55
	a8b8g8r8_sint_pack32                        = 56
	a8b8g8r8_srgb_pack32                        = 57
	a2r10g10b10_unorm_pack32                    = 58
	a2r10g10b10_snorm_pack32                    = 59
	a2r10g10b10_uscaled_pack32                  = 60
	a2r10g10b10_sscaled_pack32                  = 61
	a2r10g10b10_uint_pack32                     = 62
	a2r10g10b10_sint_pack32                     = 63
	a2b10g10r10_unorm_pack32                    = 64
	a2b10g10r10_snorm_pack32                    = 65
	a2b10g10r10_uscaled_pack32                  = 66
	a2b10g10r10_sscaled_pack32                  = 67
	a2b10g10r10_uint_pack32                     = 68
	a2b10g10r10_sint_pack32                     = 69
	r16_unorm                                   = 70
	r16_snorm                                   = 71
	r16_uscaled                                 = 72
	r16_sscaled                                 = 73
	r16_uint                                    = 74
	r16_sint                                    = 75
	r16_sfloat                                  = 76
	r16g16_unorm                                = 77
	r16g16_snorm                                = 78
	r16g16_uscaled                              = 79
	r16g16_sscaled                              = 80
	r16g16_uint                                 = 81
	r16g16_sint                                 = 82
	r16g16_sfloat                               = 83
	r16g16b16_unorm                             = 84
	r16g16b16_snorm                             = 85
	r16g16b16_uscaled                           = 86
	r16g16b16_sscaled                           = 87
	r16g16b16_uint                              = 88
	r16g16b16_sint                              = 89
	r16g16b16_sfloat                            = 90
	r16g16b16a16_unorm                          = 91
	r16g16b16a16_snorm                          = 92
	r16g16b16a16_uscaled                        = 93
	r16g16b16a16_sscaled                        = 94
	r16g16b16a16_uint                           = 95
	r16g16b16a16_sint                           = 96
	r16g16b16a16_sfloat                         = 97
	r32_uint                                    = 98
	r32_sint                                    = 99
	r32_sfloat                                  = 100
	r32g32_uint                                 = 101
	r32g32_sint                                 = 102
	r32g32_sfloat                               = 103
	r32g32b32_uint                              = 104
	r32g32b32_sint                              = 105
	r32g32b32_sfloat                            = 106
	r32g32b32a32_uint                           = 107
	r32g32b32a32_sint                           = 108
	r32g32b32a32_sfloat                         = 109
	r64_uint                                    = 110
	r64_sint                                    = 111
	r64_sfloat                                  = 112
	r64g64_uint                                 = 113
	r64g64_sint                                 = 114
	r64g64_sfloat                               = 115
	r64g64b64_uint                              = 116
	r64g64b64_sint                              = 117
	r64g64b64_sfloat                            = 118
	r64g64b64a64_uint                           = 119
	r64g64b64a64_sint                           = 120
	r64g64b64a64_sfloat                         = 121
	b10g11r11_ufloat_pack32                     = 122
	e5b9g9r9_ufloat_pack32                      = 123
	d16_unorm                                   = 124
	x8_d24_unorm_pack32                         = 125
	d32_sfloat                                  = 126
	s8_uint                                     = 127
	d16_unorm_s8_uint                           = 128
	d24_unorm_s8_uint                           = 129
	d32_sfloat_s8_uint                          = 130
	bc1_rgb_unorm_block                         = 131
	bc1_rgb_srgb_block                          = 132
	bc1_rgba_unorm_block                        = 133
	bc1_rgba_srgb_block                         = 134
	bc2_unorm_block                             = 135
	bc2_srgb_block                              = 136
	bc3_unorm_block                             = 137
	bc3_srgb_block                              = 138
	bc4_unorm_block                             = 139
	bc4_snorm_block                             = 140
	bc5_unorm_block                             = 141
	bc5_snorm_block                             = 142
	bc6h_ufloat_block                           = 143
	bc6h_sfloat_block                           = 144
	bc7_unorm_block                             = 145
	bc7_srgb_block                              = 146
	etc2_r8g8b8_unorm_block                     = 147
	etc2_r8g8b8_srgb_block                      = 148
	etc2_r8g8b8a1_unorm_block                   = 149
	etc2_r8g8b8a1_srgb_block                    = 150
	etc2_r8g8b8a8_unorm_block                   = 151
	etc2_r8g8b8a8_srgb_block                    = 152
	eac_r11_unorm_block                         = 153
	eac_r11_snorm_block                         = 154
	eac_r11g11_unorm_block                      = 155
	eac_r11g11_snorm_block                      = 156
	astc4x4_unorm_block                         = 157
	astc4x4_srgb_block                          = 158
	astc5x4_unorm_block                         = 159
	astc5x4_srgb_block                          = 160
	astc5x5_unorm_block                         = 161
	astc5x5_srgb_block                          = 162
	astc6x5_unorm_block                         = 163
	astc6x5_srgb_block                          = 164
	astc6x6_unorm_block                         = 165
	astc6x6_srgb_block                          = 166
	astc8x5_unorm_block                         = 167
	astc8x5_srgb_block                          = 168
	astc8x6_unorm_block                         = 169
	astc8x6_srgb_block                          = 170
	astc8x8_unorm_block                         = 171
	astc8x8_srgb_block                          = 172
	astc10x5_unorm_block                        = 173
	astc10x5_srgb_block                         = 174
	astc10x6_unorm_block                        = 175
	astc10x6_srgb_block                         = 176
	astc10x8_unorm_block                        = 177
	astc10x8_srgb_block                         = 178
	astc10x10_unorm_block                       = 179
	astc10x10_srgb_block                        = 180
	astc12x10_unorm_block                       = 181
	astc12x10_srgb_block                        = 182
	astc12x12_unorm_block                       = 183
	astc12x12_srgb_block                        = 184
	g8b8g8r8_422_unorm                          = 1000156000
	b8g8r8g8_422_unorm                          = 1000156001
	g8_b8_r8_3plane420_unorm                    = 1000156002
	g8_b8r8_2plane420_unorm                     = 1000156003
	g8_b8_r8_3plane422_unorm                    = 1000156004
	g8_b8r8_2plane422_unorm                     = 1000156005
	g8_b8_r8_3plane444_unorm                    = 1000156006
	r10x6_unorm_pack16                          = 1000156007
	r10x6g10x6_unorm2pack16                     = 1000156008
	r10x6g10x6b10x6a10x6_unorm4pack16           = 1000156009
	g10x6b10x6g10x6r10x6_422_unorm4pack16       = 1000156010
	b10x6g10x6r10x6g10x6_422_unorm4pack16       = 1000156011
	g10x6_b10x6_r10x6_3plane420_unorm3pack16    = 1000156012
	g10x6_b10x6r10x6_2plane420_unorm3pack16     = 1000156013
	g10x6_b10x6_r10x6_3plane422_unorm3pack16    = 1000156014
	g10x6_b10x6r10x6_2plane422_unorm3pack16     = 1000156015
	g10x6_b10x6_r10x6_3plane444_unorm3pack16    = 1000156016
	r12x4_unorm_pack16                          = 1000156017
	r12x4g12x4_unorm2pack16                     = 1000156018
	r12x4g12x4b12x4a12x4_unorm4pack16           = 1000156019
	g12x4b12x4g12x4r12x4_422_unorm4pack16       = 1000156020
	b12x4g12x4r12x4g12x4_422_unorm4pack16       = 1000156021
	g12x4_b12x4_r12x4_3plane420_unorm3pack16    = 1000156022
	g12x4_b12x4r12x4_2plane420_unorm3pack16     = 1000156023
	g12x4_b12x4_r12x4_3plane422_unorm3pack16    = 1000156024
	g12x4_b12x4r12x4_2plane422_unorm3pack16     = 1000156025
	g12x4_b12x4_r12x4_3plane444_unorm3pack16    = 1000156026
	g16b16g16r16_422_unorm                      = 1000156027
	b16g16r16g16_422_unorm                      = 1000156028
	g16_b16_r16_3plane420_unorm                 = 1000156029
	g16_b16r16_2plane420_unorm                  = 1000156030
	g16_b16_r16_3plane422_unorm                 = 1000156031
	g16_b16r16_2plane422_unorm                  = 1000156032
	g16_b16_r16_3plane444_unorm                 = 1000156033
	g8_b8r8_2plane444_unorm                     = 1000330000
	g10x6_b10x6r10x6_2plane444_unorm3pack16     = 1000330001
	g12x4_b12x4r12x4_2plane444_unorm3pack16     = 1000330002
	g16_b16r16_2plane444_unorm                  = 1000330003
	a4r4g4b4_unorm_pack16                       = 1000340000
	a4b4g4r4_unorm_pack16                       = 1000340001
	astc4x4_sfloat_block                        = 1000066000
	astc5x4_sfloat_block                        = 1000066001
	astc5x5_sfloat_block                        = 1000066002
	astc6x5_sfloat_block                        = 1000066003
	astc6x6_sfloat_block                        = 1000066004
	astc8x5_sfloat_block                        = 1000066005
	astc8x6_sfloat_block                        = 1000066006
	astc8x8_sfloat_block                        = 1000066007
	astc10x5_sfloat_block                       = 1000066008
	astc10x6_sfloat_block                       = 1000066009
	astc10x8_sfloat_block                       = 1000066010
	astc10x10_sfloat_block                      = 1000066011
	astc12x10_sfloat_block                      = 1000066012
	astc12x12_sfloat_block                      = 1000066013
	a1b5g5r5_unorm_pack16                       = 1000470000
	a8_unorm                                    = 1000470001
	pvrtc1_2bpp_unorm_block_img                 = 1000054000
	pvrtc1_4bpp_unorm_block_img                 = 1000054001
	pvrtc2_2bpp_unorm_block_img                 = 1000054002
	pvrtc2_4bpp_unorm_block_img                 = 1000054003
	pvrtc1_2bpp_srgb_block_img                  = 1000054004
	pvrtc1_4bpp_srgb_block_img                  = 1000054005
	pvrtc2_2bpp_srgb_block_img                  = 1000054006
	pvrtc2_4bpp_srgb_block_img                  = 1000054007
	r8_bool_arm                                 = 1000460000
	r16g16_sfixed5_nv                           = 1000464000
	r10x6_uint_pack16_arm                       = 1000609000
	r10x6g10x6_uint2pack16_arm                  = 1000609001
	r10x6g10x6b10x6a10x6_uint4pack16_arm        = 1000609002
	r12x4_uint_pack16_arm                       = 1000609003
	r12x4g12x4_uint2pack16_arm                  = 1000609004
	r12x4g12x4b12x4a12x4_uint4pack16_arm        = 1000609005
	r14x2_uint_pack16_arm                       = 1000609006
	r14x2g14x2_uint2pack16_arm                  = 1000609007
	r14x2g14x2b14x2a14x2_uint4pack16_arm        = 1000609008
	r14x2_unorm_pack16_arm                      = 1000609009
	r14x2g14x2_unorm2pack16_arm                 = 1000609010
	r14x2g14x2b14x2a14x2_unorm4pack16_arm       = 1000609011
	g14x2_b14x2r14x2_2plane420_unorm3pack16_arm = 1000609012
	g14x2_b14x2r14x2_2plane422_unorm3pack16_arm = 1000609013
	max_enum                                    = max_int
}

pub enum ImageTiling as u32 {
	optimal                 = 0
	linear                  = 1
	drm_format_modifier_ext = 1000158000
	max_enum                = max_int
}

pub enum ImageType as u32 {
	_1d      = 0
	_2d      = 1
	_3d      = 2
	max_enum = max_int
}

pub enum PhysicalDeviceType as u32 {
	other          = 0
	integrated_gpu = 1
	discrete_gpu   = 2
	virtual_gpu    = 3
	cpu            = 4
	max_enum       = max_int
}

pub enum QueryType as u32 {
	occlusion                                                      = 0
	pipeline_statistics                                            = 1
	timestamp                                                      = 2
	result_status_only_khr                                         = 1000023000
	transform_feedback_stream_ext                                  = 1000028004
	performance_query_khr                                          = 1000116000
	acceleration_structure_compacted_size_khr                      = 1000150000
	acceleration_structure_serialization_size_khr                  = 1000150001
	acceleration_structure_compacted_size_nv                       = 1000165000
	performance_query_intel                                        = 1000210000
	video_encode_feedback_khr                                      = 1000299000
	mesh_primitives_generated_ext                                  = 1000328000
	primitives_generated_ext                                       = 1000382000
	acceleration_structure_serialization_bottom_level_pointers_khr = 1000386000
	acceleration_structure_size_khr                                = 1000386001
	micromap_serialization_size_ext                                = 1000396000
	micromap_compacted_size_ext                                    = 1000396001
	max_enum                                                       = max_int
}

pub enum SharingMode as u32 {
	exclusive  = 0
	concurrent = 1
	max_enum   = max_int
}

pub enum ComponentSwizzle as u32 {
	identity = 0
	zero     = 1
	one      = 2
	r        = 3
	g        = 4
	b        = 5
	a        = 6
	max_enum = max_int
}

pub enum ImageViewType as u32 {
	_1d        = 0
	_2d        = 1
	_3d        = 2
	cube       = 3
	_1d_array  = 4
	_2d_array  = 5
	cube_array = 6
	max_enum   = max_int
}

pub enum CommandBufferLevel as u32 {
	primary   = 0
	secondary = 1
	max_enum  = max_int
}

pub enum IndexType as u32 {
	uint16   = 0
	uint32   = 1
	uint8    = 1000265000
	none_khr = 1000165000
	max_enum = max_int
}

pub enum PipelineCacheHeaderVersion as u32 {
	one      = 1
	max_enum = max_int
}

pub enum BorderColor as u32 {
	float_transparent_black = 0
	int_transparent_black   = 1
	float_opaque_black      = 2
	int_opaque_black        = 3
	float_opaque_white      = 4
	int_opaque_white        = 5
	float_custom_ext        = 1000287003
	int_custom_ext          = 1000287004
	max_enum                = max_int
}

pub enum Filter as u32 {
	nearest   = 0
	linear    = 1
	cubic_ext = 1000015000
	max_enum  = max_int
}

pub enum SamplerAddressMode as u32 {
	repeat               = 0
	mirrored_repeat      = 1
	clamp_to_edge        = 2
	clamp_to_border      = 3
	mirror_clamp_to_edge = 4
	max_enum             = max_int
}

pub enum SamplerMipmapMode as u32 {
	nearest  = 0
	linear   = 1
	max_enum = max_int
}

pub enum CompareOp as u32 {
	never            = 0
	less             = 1
	equal            = 2
	less_or_equal    = 3
	greater          = 4
	not_equal        = 5
	greater_or_equal = 6
	always           = 7
	max_enum         = max_int
}

pub enum DescriptorType as u32 {
	sampler                               = 0
	combined_image_sampler                = 1
	sampled_image                         = 2
	storage_image                         = 3
	uniform_texel_buffer                  = 4
	storage_texel_buffer                  = 5
	uniform_buffer                        = 6
	storage_buffer                        = 7
	uniform_buffer_dynamic                = 8
	storage_buffer_dynamic                = 9
	input_attachment                      = 10
	inline_uniform_block                  = 1000138000
	acceleration_structure_khr            = 1000150000
	acceleration_structure_nv             = 1000165000
	sample_weight_image_qcom              = 1000440000
	block_match_image_qcom                = 1000440001
	tensor_arm                            = 1000460000
	mutable_ext                           = 1000351000
	partitioned_acceleration_structure_nv = 1000570000
	max_enum                              = max_int
}

pub enum PipelineBindPoint as u32 {
	graphics               = 0
	compute                = 1
	ray_tracing_khr        = 1000165000
	subpass_shading_huawei = 1000369003
	data_graph_arm         = 1000507000
	max_enum               = max_int
}

pub enum BlendFactor as u32 {
	zero                     = 0
	one                      = 1
	src_color                = 2
	one_minus_src_color      = 3
	dst_color                = 4
	one_minus_dst_color      = 5
	src_alpha                = 6
	one_minus_src_alpha      = 7
	dst_alpha                = 8
	one_minus_dst_alpha      = 9
	constant_color           = 10
	one_minus_constant_color = 11
	constant_alpha           = 12
	one_minus_constant_alpha = 13
	src_alpha_saturate       = 14
	src1_color               = 15
	one_minus_src1_color     = 16
	src1_alpha               = 17
	one_minus_src1_alpha     = 18
	max_enum                 = max_int
}

pub enum BlendOp as u32 {
	add                    = 0
	subtract               = 1
	reverse_subtract       = 2
	min                    = 3
	max                    = 4
	zero_ext               = 1000148000
	src_ext                = 1000148001
	dst_ext                = 1000148002
	src_over_ext           = 1000148003
	dst_over_ext           = 1000148004
	src_in_ext             = 1000148005
	dst_in_ext             = 1000148006
	src_out_ext            = 1000148007
	dst_out_ext            = 1000148008
	src_atop_ext           = 1000148009
	dst_atop_ext           = 1000148010
	xor_ext                = 1000148011
	multiply_ext           = 1000148012
	screen_ext             = 1000148013
	overlay_ext            = 1000148014
	darken_ext             = 1000148015
	lighten_ext            = 1000148016
	colordodge_ext         = 1000148017
	colorburn_ext          = 1000148018
	hardlight_ext          = 1000148019
	softlight_ext          = 1000148020
	difference_ext         = 1000148021
	exclusion_ext          = 1000148022
	invert_ext             = 1000148023
	invert_rgb_ext         = 1000148024
	lineardodge_ext        = 1000148025
	linearburn_ext         = 1000148026
	vividlight_ext         = 1000148027
	linearlight_ext        = 1000148028
	pinlight_ext           = 1000148029
	hardmix_ext            = 1000148030
	hsl_hue_ext            = 1000148031
	hsl_saturation_ext     = 1000148032
	hsl_color_ext          = 1000148033
	hsl_luminosity_ext     = 1000148034
	plus_ext               = 1000148035
	plus_clamped_ext       = 1000148036
	plus_clamped_alpha_ext = 1000148037
	plus_darker_ext        = 1000148038
	minus_ext              = 1000148039
	minus_clamped_ext      = 1000148040
	contrast_ext           = 1000148041
	invert_ovg_ext         = 1000148042
	red_ext                = 1000148043
	green_ext              = 1000148044
	blue_ext               = 1000148045
	max_enum               = max_int
}

pub enum DynamicState as u32 {
	viewport                                = 0
	scissor                                 = 1
	line_width                              = 2
	depth_bias                              = 3
	blend_constants                         = 4
	depth_bounds                            = 5
	stencil_compare_mask                    = 6
	stencil_write_mask                      = 7
	stencil_reference                       = 8
	cull_mode                               = 1000267000
	front_face                              = 1000267001
	primitive_topology                      = 1000267002
	viewport_with_count                     = 1000267003
	scissor_with_count                      = 1000267004
	vertex_input_binding_stride             = 1000267005
	depth_test_enable                       = 1000267006
	depth_write_enable                      = 1000267007
	depth_compare_op                        = 1000267008
	depth_bounds_test_enable                = 1000267009
	stencil_test_enable                     = 1000267010
	stencil_op                              = 1000267011
	rasterizer_discard_enable               = 1000377001
	depth_bias_enable                       = 1000377002
	primitive_restart_enable                = 1000377004
	line_stipple                            = 1000259000
	viewport_w_scaling_nv                   = 1000087000
	discard_rectangle_ext                   = 1000099000
	discard_rectangle_enable_ext            = 1000099001
	discard_rectangle_mode_ext              = 1000099002
	sample_locations_ext                    = 1000143000
	ray_tracing_pipeline_stack_size_khr     = 1000347000
	viewport_shading_rate_palette_nv        = 1000164004
	viewport_coarse_sample_order_nv         = 1000164006
	exclusive_scissor_enable_nv             = 1000205000
	exclusive_scissor_nv                    = 1000205001
	fragment_shading_rate_khr               = 1000226000
	vertex_input_ext                        = 1000352000
	patch_control_points_ext                = 1000377000
	logic_op_ext                            = 1000377003
	color_write_enable_ext                  = 1000381000
	depth_clamp_enable_ext                  = 1000455003
	polygon_mode_ext                        = 1000455004
	rasterization_samples_ext               = 1000455005
	sample_mask_ext                         = 1000455006
	alpha_to_coverage_enable_ext            = 1000455007
	alpha_to_one_enable_ext                 = 1000455008
	logic_op_enable_ext                     = 1000455009
	color_blend_enable_ext                  = 1000455010
	color_blend_equation_ext                = 1000455011
	color_write_mask_ext                    = 1000455012
	tessellation_domain_origin_ext          = 1000455002
	rasterization_stream_ext                = 1000455013
	conservative_rasterization_mode_ext     = 1000455014
	extra_primitive_overestimation_size_ext = 1000455015
	depth_clip_enable_ext                   = 1000455016
	sample_locations_enable_ext             = 1000455017
	color_blend_advanced_ext                = 1000455018
	provoking_vertex_mode_ext               = 1000455019
	line_rasterization_mode_ext             = 1000455020
	line_stipple_enable_ext                 = 1000455021
	depth_clip_negative_one_to_one_ext      = 1000455022
	viewport_w_scaling_enable_nv            = 1000455023
	viewport_swizzle_nv                     = 1000455024
	coverage_to_color_enable_nv             = 1000455025
	coverage_to_color_location_nv           = 1000455026
	coverage_modulation_mode_nv             = 1000455027
	coverage_modulation_table_enable_nv     = 1000455028
	coverage_modulation_table_nv            = 1000455029
	shading_rate_image_enable_nv            = 1000455030
	representative_fragment_test_enable_nv  = 1000455031
	coverage_reduction_mode_nv              = 1000455032
	attachment_feedback_loop_enable_ext     = 1000524000
	depth_clamp_range_ext                   = 1000582000
	max_enum                                = max_int
}

pub enum FrontFace as u32 {
	counter_clockwise = 0
	clockwise         = 1
	max_enum          = max_int
}

pub enum VertexInputRate as u32 {
	vertex   = 0
	instance = 1
	max_enum = max_int
}

pub enum PrimitiveTopology as u32 {
	point_list                    = 0
	line_list                     = 1
	line_strip                    = 2
	triangle_list                 = 3
	triangle_strip                = 4
	triangle_fan                  = 5
	line_list_with_adjacency      = 6
	line_strip_with_adjacency     = 7
	triangle_list_with_adjacency  = 8
	triangle_strip_with_adjacency = 9
	patch_list                    = 10
	max_enum                      = max_int
}

pub enum PolygonMode as u32 {
	fill              = 0
	line              = 1
	point             = 2
	fill_rectangle_nv = 1000153000
	max_enum          = max_int
}

pub enum StencilOp as u32 {
	keep                = 0
	zero                = 1
	replace             = 2
	increment_and_clamp = 3
	decrement_and_clamp = 4
	invert              = 5
	increment_and_wrap  = 6
	decrement_and_wrap  = 7
	max_enum            = max_int
}

pub enum LogicOp as u32 {
	clear         = 0
	and           = 1
	and_reverse   = 2
	copy          = 3
	and_inverted  = 4
	no            = 5
	xor           = 6
	or            = 7
	nor           = 8
	equivalent    = 9
	invert        = 10
	or_reverse    = 11
	copy_inverted = 12
	or_inverted   = 13
	nand          = 14
	set           = 15
	max_enum      = max_int
}

pub enum AttachmentLoadOp as u32 {
	load      = 0
	clear     = 1
	dont_care = 2
	none      = 1000400000
	max_enum  = max_int
}

pub enum AttachmentStoreOp as u32 {
	store     = 0
	dont_care = 1
	none      = 1000301000
	max_enum  = max_int
}

pub enum SubpassContents as u32 {
	inline                                   = 0
	secondary_command_buffers                = 1
	inline_and_secondary_command_buffers_khr = 1000451000
	max_enum                                 = max_int
}

pub enum AccessFlagBits as u32 {
	indirect_command_read                     = u32(0x00000001)
	index_read                                = u32(0x00000002)
	vertex_attribute_read                     = u32(0x00000004)
	uniform_read                              = u32(0x00000008)
	input_attachment_read                     = u32(0x00000010)
	shader_read                               = u32(0x00000020)
	shader_write                              = u32(0x00000040)
	color_attachment_read                     = u32(0x00000080)
	color_attachment_write                    = u32(0x00000100)
	depth_stencil_attachment_read             = u32(0x00000200)
	depth_stencil_attachment_write            = u32(0x00000400)
	transfer_read                             = u32(0x00000800)
	transfer_write                            = u32(0x00001000)
	host_read                                 = u32(0x00002000)
	host_write                                = u32(0x00004000)
	memory_read                               = u32(0x00008000)
	memory_write                              = u32(0x00010000)
	none                                      = 0
	transform_feedback_write_bit_ext          = u32(0x02000000)
	transform_feedback_counter_read_bit_ext   = u32(0x04000000)
	transform_feedback_counter_write_bit_ext  = u32(0x08000000)
	conditional_rendering_read_bit_ext        = u32(0x00100000)
	color_attachment_read_noncoherent_bit_ext = u32(0x00080000)
	acceleration_structure_read               = u32(0x00200000)
	acceleration_structure_write              = u32(0x00400000)
	fragment_density_map_read_bit_ext         = u32(0x01000000)
	fragment_shading_rate_attachment_read     = u32(0x00800000)
	command_preprocess_read_bit_ext           = u32(0x00020000)
	command_preprocess_write_bit_ext          = u32(0x00040000)
	max_enum                                  = max_int
}
pub type AccessFlags = u32

pub enum ImageAspectFlagBits as u32 {
	color                 = u32(0x00000001)
	depth                 = u32(0x00000002)
	stencil               = u32(0x00000004)
	metadata              = u32(0x00000008)
	plane0                = u32(0x00000010)
	plane1                = u32(0x00000020)
	plane2                = u32(0x00000040)
	none                  = 0
	memory_plane0_bit_ext = u32(0x00000080)
	memory_plane1_bit_ext = u32(0x00000100)
	memory_plane2_bit_ext = u32(0x00000200)
	memory_plane3_bit_ext = u32(0x00000400)
	max_enum              = max_int
}
pub type ImageAspectFlags = u32

pub enum FormatFeatureFlagBits as u32 {
	sampled_image                                                           = u32(0x00000001)
	storage_image                                                           = u32(0x00000002)
	storage_image_atomic                                                    = u32(0x00000004)
	uniform_texel_buffer                                                    = u32(0x00000008)
	storage_texel_buffer                                                    = u32(0x00000010)
	storage_texel_buffer_atomic                                             = u32(0x00000020)
	vertex_buffer                                                           = u32(0x00000040)
	color_attachment                                                        = u32(0x00000080)
	color_attachment_blend                                                  = u32(0x00000100)
	depth_stencil_attachment                                                = u32(0x00000200)
	blit_src                                                                = u32(0x00000400)
	blit_dst                                                                = u32(0x00000800)
	sampled_image_filter_linear                                             = u32(0x00001000)
	transfer_src                                                            = u32(0x00004000)
	transfer_dst                                                            = u32(0x00008000)
	midpoint_chroma_samples                                                 = u32(0x00020000)
	sampled_image_ycbcr_conversion_linear_filter                            = u32(0x00040000)
	sampled_image_ycbcr_conversion_separate_reconstruction_filter           = u32(0x00080000)
	sampled_image_ycbcr_conversion_chroma_reconstruction_explicit           = u32(0x00100000)
	sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_forceable = u32(0x00200000)
	disjoint                                                                = u32(0x00400000)
	cosited_chroma_samples                                                  = u32(0x00800000)
	sampled_image_filter_minmax                                             = u32(0x00010000)
	video_decode_output                                                     = u32(0x02000000)
	video_decode_dpb                                                        = u32(0x04000000)
	acceleration_structure_vertex_buffer                                    = u32(0x20000000)
	sampled_image_filter_cubic_bit_ext                                      = u32(0x00002000)
	fragment_density_map_bit_ext                                            = u32(0x01000000)
	fragment_shading_rate_attachment                                        = u32(0x40000000)
	video_encode_input                                                      = u32(0x08000000)
	video_encode_dpb                                                        = u32(0x10000000)
	max_enum                                                                = max_int
}
pub type FormatFeatureFlags = u32

pub enum ImageCreateFlagBits as u32 {
	sparse_binding                                = u32(0x00000001)
	sparse_residency                              = u32(0x00000002)
	sparse_aliased                                = u32(0x00000004)
	mutable_format                                = u32(0x00000008)
	cube_compatible                               = u32(0x00000010)
	alias                                         = u32(0x00000400)
	split_instance_bind_regions                   = u32(0x00000040)
	_2d_array_compatible                          = u32(0x00000020)
	block_texel_view_compatible                   = u32(0x00000080)
	extended_usage                                = u32(0x00000100)
	protected                                     = u32(0x00000800)
	disjoint                                      = u32(0x00000200)
	corner_sampled_bit_nv                         = u32(0x00002000)
	sample_locations_compatible_depth_bit_ext     = u32(0x00001000)
	subsampled_bit_ext                            = u32(0x00004000)
	descriptor_buffer_capture_replay_bit_ext      = u32(0x00010000)
	multisampled_render_to_single_sampled_bit_ext = u32(0x00040000)
	_2d_view_compatible_bit_ext                   = u32(0x00020000)
	video_profile_independent                     = u32(0x00100000)
	fragment_density_map_offset_bit_ext           = u32(0x00008000)
	max_enum                                      = max_int
}
pub type ImageCreateFlags = u32

pub enum SampleCountFlagBits as u32 {
	_1       = u32(0x00000001)
	_2       = u32(0x00000002)
	_4       = u32(0x00000004)
	_8       = u32(0x00000008)
	_16      = u32(0x00000010)
	_32      = u32(0x00000020)
	_64      = u32(0x00000040)
	max_enum = max_int
}
pub type SampleCountFlags = u32

pub enum ImageUsageFlagBits as u32 {
	transfer_src                        = u32(0x00000001)
	transfer_dst                        = u32(0x00000002)
	sampled                             = u32(0x00000004)
	storage                             = u32(0x00000008)
	color_attachment                    = u32(0x00000010)
	depth_stencil_attachment            = u32(0x00000020)
	transient_attachment                = u32(0x00000040)
	input_attachment                    = u32(0x00000080)
	host_transfer                       = u32(0x00400000)
	video_decode_dst                    = u32(0x00000400)
	video_decode_src                    = u32(0x00000800)
	video_decode_dpb                    = u32(0x00001000)
	fragment_density_map_bit_ext        = u32(0x00000200)
	fragment_shading_rate_attachment    = u32(0x00000100)
	video_encode_dst                    = u32(0x00002000)
	video_encode_src                    = u32(0x00004000)
	video_encode_dpb                    = u32(0x00008000)
	attachment_feedback_loop_bit_ext    = u32(0x00080000)
	invocation_mask_bit_huawei          = u32(0x00040000)
	sample_weight_bit_qcom              = u32(0x00100000)
	sample_block_match_bit_qcom         = u32(0x00200000)
	tensor_aliasing_bit_arm             = u32(0x00800000)
	tile_memory_bit_qcom                = u32(0x08000000)
	video_encode_quantization_delta_map = u32(0x02000000)
	video_encode_emphasis_map           = u32(0x04000000)
	max_enum                            = max_int
}
pub type ImageUsageFlags = u32

pub enum InstanceCreateFlagBits as u32 {
	enumerate_portability = u32(0x00000001)
	max_enum              = max_int
}
pub type InstanceCreateFlags = u32

pub enum MemoryHeapFlagBits as u32 {
	device_local         = u32(0x00000001)
	multi_instance       = u32(0x00000002)
	tile_memory_bit_qcom = u32(0x00000008)
	max_enum             = max_int
}
pub type MemoryHeapFlags = u32

pub enum MemoryPropertyFlagBits as u32 {
	device_local            = u32(0x00000001)
	host_visible            = u32(0x00000002)
	host_coherent           = u32(0x00000004)
	host_cached             = u32(0x00000008)
	lazily_allocated        = u32(0x00000010)
	protected               = u32(0x00000020)
	device_coherent_bit_amd = u32(0x00000040)
	device_uncached_bit_amd = u32(0x00000080)
	rdma_capable_bit_nv     = u32(0x00000100)
	max_enum                = max_int
}
pub type MemoryPropertyFlags = u32

pub enum QueueFlagBits as u32 {
	graphics            = u32(0x00000001)
	compute             = u32(0x00000002)
	transfer            = u32(0x00000004)
	sparse_binding      = u32(0x00000008)
	protected           = u32(0x00000010)
	video_decode        = u32(0x00000020)
	video_encode        = u32(0x00000040)
	optical_flow_bit_nv = u32(0x00000100)
	data_graph_bit_arm  = u32(0x00000400)
	max_enum            = max_int
}
pub type QueueFlags = u32
pub type DeviceCreateFlags = u32

pub enum DeviceQueueCreateFlagBits as u32 {
	protected = u32(0x00000001)
	max_enum  = max_int
}
pub type DeviceQueueCreateFlags = u32

pub enum PipelineStageFlagBits as u32 {
	top_of_pipe                      = u32(0x00000001)
	draw_indirect                    = u32(0x00000002)
	vertex_input                     = u32(0x00000004)
	vertex_shader                    = u32(0x00000008)
	tessellation_control_shader      = u32(0x00000010)
	tessellation_evaluation_shader   = u32(0x00000020)
	geometry_shader                  = u32(0x00000040)
	fragment_shader                  = u32(0x00000080)
	early_fragment_tests             = u32(0x00000100)
	late_fragment_tests              = u32(0x00000200)
	color_attachment_output          = u32(0x00000400)
	compute_shader                   = u32(0x00000800)
	transfer                         = u32(0x00001000)
	bottom_of_pipe                   = u32(0x00002000)
	host                             = u32(0x00004000)
	all_graphics                     = u32(0x00008000)
	all_commands                     = u32(0x00010000)
	none                             = 0
	transform_feedback_bit_ext       = u32(0x01000000)
	conditional_rendering_bit_ext    = u32(0x00040000)
	acceleration_structure_build     = u32(0x02000000)
	ray_tracing_shader               = u32(0x00200000)
	fragment_density_process_bit_ext = u32(0x00800000)
	fragment_shading_rate_attachment = u32(0x00400000)
	task_shader_bit_ext              = u32(0x00080000)
	mesh_shader_bit_ext              = u32(0x00100000)
	command_preprocess_bit_ext       = u32(0x00020000)
	max_enum                         = max_int
}
pub type PipelineStageFlags = u32

pub enum MemoryMapFlagBits as u32 {
	placed_bit_ext = u32(0x00000001)
	max_enum       = max_int
}
pub type MemoryMapFlags = u32

pub enum SparseMemoryBindFlagBits as u32 {
	metadata = u32(0x00000001)
	max_enum = max_int
}
pub type SparseMemoryBindFlags = u32

pub enum SparseImageFormatFlagBits as u32 {
	single_miptail         = u32(0x00000001)
	aligned_mip_size       = u32(0x00000002)
	nonstandard_block_size = u32(0x00000004)
	max_enum               = max_int
}
pub type SparseImageFormatFlags = u32

pub enum FenceCreateFlagBits as u32 {
	signaled = u32(0x00000001)
	max_enum = max_int
}
pub type FenceCreateFlags = u32
pub type SemaphoreCreateFlags = u32

pub enum QueryPoolCreateFlagBits as u32 {
	reset    = u32(0x00000001)
	max_enum = max_int
}
pub type QueryPoolCreateFlags = u32

pub enum QueryPipelineStatisticFlagBits as u32 {
	input_assembly_vertices                       = u32(0x00000001)
	input_assembly_primitives                     = u32(0x00000002)
	vertex_shader_invocations                     = u32(0x00000004)
	geometry_shader_invocations                   = u32(0x00000008)
	geometry_shader_primitives                    = u32(0x00000010)
	clipping_invocations                          = u32(0x00000020)
	clipping_primitives                           = u32(0x00000040)
	fragment_shader_invocations                   = u32(0x00000080)
	tessellation_control_shader_patches           = u32(0x00000100)
	tessellation_evaluation_shader_invocations    = u32(0x00000200)
	compute_shader_invocations                    = u32(0x00000400)
	task_shader_invocations_bit_ext               = u32(0x00000800)
	mesh_shader_invocations_bit_ext               = u32(0x00001000)
	cluster_culling_shader_invocations_bit_huawei = u32(0x00002000)
	max_enum                                      = max_int
}
pub type QueryPipelineStatisticFlags = u32

pub enum QueryResultFlagBits as u32 {
	_64               = u32(0x00000001)
	wait              = u32(0x00000002)
	with_availability = u32(0x00000004)
	partial           = u32(0x00000008)
	with_status       = u32(0x00000010)
	max_enum          = max_int
}
pub type QueryResultFlags = u32

pub enum BufferCreateFlagBits as u32 {
	sparse_binding                           = u32(0x00000001)
	sparse_residency                         = u32(0x00000002)
	sparse_aliased                           = u32(0x00000004)
	protected                                = u32(0x00000008)
	device_address_capture_replay            = u32(0x00000010)
	descriptor_buffer_capture_replay_bit_ext = u32(0x00000020)
	video_profile_independent                = u32(0x00000040)
	max_enum                                 = max_int
}
pub type BufferCreateFlags = u32

pub enum BufferUsageFlagBits as u32 {
	transfer_src                                 = u32(0x00000001)
	transfer_dst                                 = u32(0x00000002)
	uniform_texel_buffer                         = u32(0x00000004)
	storage_texel_buffer                         = u32(0x00000008)
	uniform_buffer                               = u32(0x00000010)
	storage_buffer                               = u32(0x00000020)
	index_buffer                                 = u32(0x00000040)
	vertex_buffer                                = u32(0x00000080)
	indirect_buffer                              = u32(0x00000100)
	shader_device_address                        = u32(0x00020000)
	video_decode_src                             = u32(0x00002000)
	video_decode_dst                             = u32(0x00004000)
	transform_feedback_buffer_bit_ext            = u32(0x00000800)
	transform_feedback_counter_buffer_bit_ext    = u32(0x00001000)
	conditional_rendering_bit_ext                = u32(0x00000200)
	acceleration_structure_build_input_read_only = u32(0x00080000)
	acceleration_structure_storage               = u32(0x00100000)
	shader_binding_table                         = u32(0x00000400)
	video_encode_dst                             = u32(0x00008000)
	video_encode_src                             = u32(0x00010000)
	sampler_descriptor_buffer_bit_ext            = u32(0x00200000)
	resource_descriptor_buffer_bit_ext           = u32(0x00400000)
	push_descriptors_descriptor_buffer_bit_ext   = u32(0x04000000)
	micromap_build_input_read_only_bit_ext       = u32(0x00800000)
	micromap_storage_bit_ext                     = u32(0x01000000)
	tile_memory_bit_qcom                         = u32(0x08000000)
	max_enum                                     = max_int
}
pub type BufferUsageFlags = u32

pub enum ImageViewCreateFlagBits as u32 {
	fragment_density_map_dynamic_bit_ext     = u32(0x00000001)
	descriptor_buffer_capture_replay_bit_ext = u32(0x00000004)
	fragment_density_map_deferred_bit_ext    = u32(0x00000002)
	max_enum                                 = max_int
}
pub type ImageViewCreateFlags = u32

pub enum DependencyFlagBits as u32 {
	by_region                                      = u32(0x00000001)
	device_group                                   = u32(0x00000004)
	view_local                                     = u32(0x00000002)
	feedback_loop_bit_ext                          = u32(0x00000008)
	queue_family_ownership_transfer_use_all_stages = u32(0x00000020)
	asymmetric_event                               = u32(0x00000040)
	max_enum                                       = max_int
}
pub type DependencyFlags = u32

pub enum CommandPoolCreateFlagBits as u32 {
	transient            = u32(0x00000001)
	reset_command_buffer = u32(0x00000002)
	protected            = u32(0x00000004)
	max_enum             = max_int
}
pub type CommandPoolCreateFlags = u32

pub enum CommandPoolResetFlagBits as u32 {
	release_resources = u32(0x00000001)
	max_enum          = max_int
}
pub type CommandPoolResetFlags = u32

pub enum CommandBufferUsageFlagBits as u32 {
	one_time_submit      = u32(0x00000001)
	render_pass_continue = u32(0x00000002)
	simultaneous_use     = u32(0x00000004)
	max_enum             = max_int
}
pub type CommandBufferUsageFlags = u32

pub enum QueryControlFlagBits as u32 {
	precise  = u32(0x00000001)
	max_enum = max_int
}
pub type QueryControlFlags = u32

pub enum CommandBufferResetFlagBits as u32 {
	release_resources = u32(0x00000001)
	max_enum          = max_int
}
pub type CommandBufferResetFlags = u32

pub enum EventCreateFlagBits as u32 {
	device_only = u32(0x00000001)
	max_enum    = max_int
}
pub type EventCreateFlags = u32
pub type BufferViewCreateFlags = u32
pub type ShaderModuleCreateFlags = u32

pub enum PipelineCacheCreateFlagBits as u32 {
	externally_synchronized       = u32(0x00000001)
	internally_synchronized_merge = u32(0x00000008)
	max_enum                      = max_int
}
pub type PipelineCacheCreateFlags = u32

pub enum PipelineCreateFlagBits as u32 {
	disable_optimization                              = u32(0x00000001)
	allow_derivatives                                 = u32(0x00000002)
	derivative                                        = u32(0x00000004)
	dispatch_base                                     = u32(0x00000010)
	view_index_from_device_index                      = u32(0x00000008)
	fail_on_pipeline_compile_required                 = u32(0x00000100)
	early_return_on_failure                           = u32(0x00000200)
	no_protected_access                               = u32(0x08000000)
	protected_access_only                             = u32(0x40000000)
	ray_tracing_no_null_any_hit_shaders               = u32(0x00004000)
	ray_tracing_no_null_closest_hit_shaders           = u32(0x00008000)
	ray_tracing_no_null_miss_shaders                  = u32(0x00010000)
	ray_tracing_no_null_intersection_shaders          = u32(0x00020000)
	ray_tracing_skip_triangles                        = u32(0x00001000)
	ray_tracing_skip_aabbs                            = u32(0x00002000)
	ray_tracing_shader_group_handle_capture_replay    = u32(0x00080000)
	defer_compile_bit_nv                              = u32(0x00000020)
	rendering_fragment_density_map_attachment_bit_ext = u32(0x00400000)
	rendering_fragment_shading_rate_attachment        = u32(0x00200000)
	capture_statistics                                = u32(0x00000040)
	capture_internal_representations                  = u32(0x00000080)
	indirect_bindable_bit_nv                          = u32(0x00040000)
	library                                           = u32(0x00000800)
	descriptor_buffer_bit_ext                         = u32(0x20000000)
	retain_link_time_optimization_info_bit_ext        = u32(0x00800000)
	link_time_optimization_bit_ext                    = u32(0x00000400)
	ray_tracing_allow_motion_bit_nv                   = u32(0x00100000)
	color_attachment_feedback_loop_bit_ext            = u32(0x02000000)
	depth_stencil_attachment_feedback_loop_bit_ext    = u32(0x04000000)
	ray_tracing_opacity_micromap_bit_ext              = u32(0x01000000)
	max_enum                                          = max_int
}
pub type PipelineCreateFlags = u32

pub enum PipelineShaderStageCreateFlagBits as u32 {
	allow_varying_subgroup_size = u32(0x00000001)
	require_full_subgroups      = u32(0x00000002)
	max_enum                    = max_int
}
pub type PipelineShaderStageCreateFlags = u32

pub enum ShaderStageFlagBits as u32 {
	vertex                     = u32(0x00000001)
	tessellation_control       = u32(0x00000002)
	tessellation_evaluation    = u32(0x00000004)
	geometry                   = u32(0x00000008)
	fragment                   = u32(0x00000010)
	compute                    = u32(0x00000020)
	all_graphics               = u32(0x0000001F)
	all                        = u32(0x7FFFFFFF)
	raygen                     = u32(0x00000100)
	any_hit                    = u32(0x00000200)
	closest_hit                = u32(0x00000400)
	miss                       = u32(0x00000800)
	intersection               = u32(0x00001000)
	callable                   = u32(0x00002000)
	task_bit_ext               = u32(0x00000040)
	mesh_bit_ext               = u32(0x00000080)
	subpass_shading_bit_huawei = u32(0x00004000)
	cluster_culling_bit_huawei = u32(0x00080000)
}

pub enum PipelineLayoutCreateFlagBits as u32 {
	independent_sets_bit_ext = u32(0x00000002)
	max_enum                 = max_int
}
pub type PipelineLayoutCreateFlags = u32
pub type ShaderStageFlags = u32

pub enum SamplerCreateFlagBits as u32 {
	subsampled_bit_ext                       = u32(0x00000001)
	subsampled_coarse_reconstruction_bit_ext = u32(0x00000002)
	descriptor_buffer_capture_replay_bit_ext = u32(0x00000008)
	non_seamless_cube_map_bit_ext            = u32(0x00000004)
	image_processing_bit_qcom                = u32(0x00000010)
	max_enum                                 = max_int
}
pub type SamplerCreateFlags = u32

pub enum DescriptorPoolCreateFlagBits as u32 {
	free_descriptor_set               = u32(0x00000001)
	update_after_bind                 = u32(0x00000002)
	host_only_bit_ext                 = u32(0x00000004)
	allow_overallocation_sets_bit_nv  = u32(0x00000008)
	allow_overallocation_pools_bit_nv = u32(0x00000010)
	max_enum                          = max_int
}
pub type DescriptorPoolCreateFlags = u32
pub type DescriptorPoolResetFlags = u32

pub enum DescriptorSetLayoutCreateFlagBits as u32 {
	update_after_bind_pool              = u32(0x00000002)
	push_descriptor                     = u32(0x00000001)
	descriptor_buffer_bit_ext           = u32(0x00000010)
	embedded_immutable_samplers_bit_ext = u32(0x00000020)
	indirect_bindable_bit_nv            = u32(0x00000080)
	host_only_pool_bit_ext              = u32(0x00000004)
	per_stage_bit_nv                    = u32(0x00000040)
	max_enum                            = max_int
}
pub type DescriptorSetLayoutCreateFlags = u32

pub enum ColorComponentFlagBits as u32 {
	r        = u32(0x00000001)
	g        = u32(0x00000002)
	b        = u32(0x00000004)
	a        = u32(0x00000008)
	max_enum = max_int
}
pub type ColorComponentFlags = u32

pub enum CullModeFlagBits as u32 {
	none           = 0
	front          = u32(0x00000001)
	back           = u32(0x00000002)
	front_and_back = u32(0x00000003)
	max_enum       = max_int
}
pub type CullModeFlags = u32
pub type PipelineVertexInputStateCreateFlags = u32
pub type PipelineInputAssemblyStateCreateFlags = u32
pub type PipelineTessellationStateCreateFlags = u32
pub type PipelineViewportStateCreateFlags = u32
pub type PipelineRasterizationStateCreateFlags = u32
pub type PipelineMultisampleStateCreateFlags = u32

pub enum PipelineDepthStencilStateCreateFlagBits as u32 {
	rasterization_order_attachment_depth_access_bit_ext   = u32(0x00000001)
	rasterization_order_attachment_stencil_access_bit_ext = u32(0x00000002)
	max_enum                                              = max_int
}
pub type PipelineDepthStencilStateCreateFlags = u32

pub enum PipelineColorBlendStateCreateFlagBits as u32 {
	rasterization_order_attachment_access_bit_ext = u32(0x00000001)
	max_enum                                      = max_int
}
pub type PipelineColorBlendStateCreateFlags = u32
pub type PipelineDynamicStateCreateFlags = u32

pub enum AttachmentDescriptionFlagBits as u32 {
	may_alias                        = u32(0x00000001)
	resolve_skip_transfer_function   = u32(0x00000002)
	resolve_enable_transfer_function = u32(0x00000004)
	max_enum                         = max_int
}
pub type AttachmentDescriptionFlags = u32

pub enum FramebufferCreateFlagBits as u32 {
	imageless = u32(0x00000001)
	max_enum  = max_int
}
pub type FramebufferCreateFlags = u32

pub enum RenderPassCreateFlagBits as u32 {
	transform_bit_qcom                   = u32(0x00000002)
	per_layer_fragment_density_bit_valve = u32(0x00000004)
	max_enum                             = max_int
}
pub type RenderPassCreateFlags = u32

pub enum SubpassDescriptionFlagBits as u32 {
	per_view_attributes_bit_nvx                           = u32(0x00000001)
	per_view_position_x_only_bit_nvx                      = u32(0x00000002)
	fragment_region_bit_qcom                              = u32(0x00000004)
	shader_resolve_bit_qcom                               = u32(0x00000008)
	tile_shading_apron_bit_qcom                           = u32(0x00000100)
	rasterization_order_attachment_color_access_bit_ext   = u32(0x00000010)
	rasterization_order_attachment_depth_access_bit_ext   = u32(0x00000020)
	rasterization_order_attachment_stencil_access_bit_ext = u32(0x00000040)
	enable_legacy_dithering_bit_ext                       = u32(0x00000080)
	max_enum                                              = max_int
}
pub type SubpassDescriptionFlags = u32

pub enum StencilFaceFlagBits as u32 {
	front          = u32(0x00000001)
	back           = u32(0x00000002)
	front_and_back = u32(0x00000003)
	max_enum       = max_int
}
pub type StencilFaceFlags = u32
pub type Extent2D = C.VkExtent2D

@[typedef]
pub struct C.VkExtent2D {
pub mut:
	width  u32
	height u32
}

pub type Extent3D = C.VkExtent3D

@[typedef]
pub struct C.VkExtent3D {
pub mut:
	width  u32
	height u32
	depth  u32
}

pub type Offset2D = C.VkOffset2D

@[typedef]
pub struct C.VkOffset2D {
pub mut:
	x i32
	y i32
}

pub type Offset3D = C.VkOffset3D

@[typedef]
pub struct C.VkOffset3D {
pub mut:
	x i32
	y i32
	z i32
}

pub type Rect2D = C.VkRect2D

@[typedef]
pub struct C.VkRect2D {
pub mut:
	offset Offset2D
	extent Extent2D
}

pub type BaseInStructure = C.VkBaseInStructure

@[typedef]
pub struct C.VkBaseInStructure {
pub mut:
	sType StructureType
	pNext &BaseInStructure
}

pub type BaseOutStructure = C.VkBaseOutStructure

@[typedef]
pub struct C.VkBaseOutStructure {
pub mut:
	sType StructureType
	pNext &BaseOutStructure
}

pub type BufferMemoryBarrier = C.VkBufferMemoryBarrier

@[typedef]
pub struct C.VkBufferMemoryBarrier {
pub mut:
	sType               StructureType = StructureType.buffer_memory_barrier
	pNext               voidptr       = unsafe { nil }
	srcAccessMask       AccessFlags
	dstAccessMask       AccessFlags
	srcQueueFamilyIndex u32
	dstQueueFamilyIndex u32
	buffer              Buffer
	offset              DeviceSize
	size                DeviceSize
}

pub type ImageSubresourceRange = C.VkImageSubresourceRange

@[typedef]
pub struct C.VkImageSubresourceRange {
pub mut:
	aspectMask     ImageAspectFlags
	baseMipLevel   u32
	levelCount     u32
	baseArrayLayer u32
	layerCount     u32
}

pub type ImageMemoryBarrier = C.VkImageMemoryBarrier

@[typedef]
pub struct C.VkImageMemoryBarrier {
pub mut:
	sType               StructureType = StructureType.image_memory_barrier
	pNext               voidptr       = unsafe { nil }
	srcAccessMask       AccessFlags
	dstAccessMask       AccessFlags
	oldLayout           ImageLayout
	newLayout           ImageLayout
	srcQueueFamilyIndex u32
	dstQueueFamilyIndex u32
	image               Image
	subresourceRange    ImageSubresourceRange
}

pub type MemoryBarrier = C.VkMemoryBarrier

@[typedef]
pub struct C.VkMemoryBarrier {
pub mut:
	sType         StructureType = StructureType.memory_barrier
	pNext         voidptr       = unsafe { nil }
	srcAccessMask AccessFlags
	dstAccessMask AccessFlags
}

pub type PFN_vkAllocationFunction = fn (voidptr, usize, usize, SystemAllocationScope)

pub type PFN_vkFreeFunction = fn (voidptr, voidptr)

pub type PFN_vkInternalAllocationNotification = fn (voidptr, usize, InternalAllocationType, SystemAllocationScope)

pub type PFN_vkInternalFreeNotification = fn (voidptr, usize, InternalAllocationType, SystemAllocationScope)

pub type PFN_vkReallocationFunction = fn (voidptr, voidptr, usize, usize, SystemAllocationScope)

pub type PFN_vkVoidFunction = fn ()

pub type AllocationCallbacks = C.VkAllocationCallbacks

@[typedef]
pub struct C.VkAllocationCallbacks {
pub mut:
	pUserData             voidptr                              = unsafe { nil }
	pfnAllocation         PFN_vkAllocationFunction             = unsafe { nil }
	pfnReallocation       PFN_vkReallocationFunction           = unsafe { nil }
	pfnFree               PFN_vkFreeFunction                   = unsafe { nil }
	pfnInternalAllocation PFN_vkInternalAllocationNotification = unsafe { nil }
	pfnInternalFree       PFN_vkInternalFreeNotification       = unsafe { nil }
}

pub type ApplicationInfo = C.VkApplicationInfo

@[typedef]
pub struct C.VkApplicationInfo {
pub mut:
	sType              StructureType = StructureType.application_info
	pNext              voidptr       = unsafe { nil }
	pApplicationName   &char
	applicationVersion u32
	pEngineName        &char
	engineVersion      u32
	apiVersion         u32
}

pub type FormatProperties = C.VkFormatProperties

@[typedef]
pub struct C.VkFormatProperties {
pub mut:
	linearTilingFeatures  FormatFeatureFlags
	optimalTilingFeatures FormatFeatureFlags
	bufferFeatures        FormatFeatureFlags
}

pub type ImageFormatProperties = C.VkImageFormatProperties

@[typedef]
pub struct C.VkImageFormatProperties {
pub mut:
	maxExtent       Extent3D
	maxMipLevels    u32
	maxArrayLayers  u32
	sampleCounts    SampleCountFlags
	maxResourceSize DeviceSize
}

pub type InstanceCreateInfo = C.VkInstanceCreateInfo

@[typedef]
pub struct C.VkInstanceCreateInfo {
pub mut:
	sType                   StructureType = StructureType.instance_create_info
	pNext                   voidptr       = unsafe { nil }
	flags                   InstanceCreateFlags
	pApplicationInfo        &ApplicationInfo
	enabledLayerCount       u32
	ppEnabledLayerNames     &&char
	enabledExtensionCount   u32
	ppEnabledExtensionNames &&char
}

pub type MemoryHeap = C.VkMemoryHeap

@[typedef]
pub struct C.VkMemoryHeap {
pub mut:
	size  DeviceSize
	flags MemoryHeapFlags
}

pub type MemoryType = C.VkMemoryType

@[typedef]
pub struct C.VkMemoryType {
pub mut:
	propertyFlags MemoryPropertyFlags
	heapIndex     u32
}

pub type PhysicalDeviceFeatures = C.VkPhysicalDeviceFeatures

@[typedef]
pub struct C.VkPhysicalDeviceFeatures {
pub mut:
	robustBufferAccess                      Bool32
	fullDrawIndexUint32                     Bool32
	imageCubeArray                          Bool32
	independentBlend                        Bool32
	geometryShader                          Bool32
	tessellationShader                      Bool32
	sampleRateShading                       Bool32
	dualSrcBlend                            Bool32
	logicOp                                 Bool32
	multiDrawIndirect                       Bool32
	drawIndirectFirstInstance               Bool32
	depthClamp                              Bool32
	depthBiasClamp                          Bool32
	fillModeNonSolid                        Bool32
	depthBounds                             Bool32
	wideLines                               Bool32
	largePoints                             Bool32
	alphaToOne                              Bool32
	multiViewport                           Bool32
	samplerAnisotropy                       Bool32
	textureCompressionETC2                  Bool32
	textureCompressionASTC_LDR              Bool32
	textureCompressionBC                    Bool32
	occlusionQueryPrecise                   Bool32
	pipelineStatisticsQuery                 Bool32
	vertexPipelineStoresAndAtomics          Bool32
	fragmentStoresAndAtomics                Bool32
	shaderTessellationAndGeometryPointSize  Bool32
	shaderImageGatherExtended               Bool32
	shaderStorageImageExtendedFormats       Bool32
	shaderStorageImageMultisample           Bool32
	shaderStorageImageReadWithoutFormat     Bool32
	shaderStorageImageWriteWithoutFormat    Bool32
	shaderUniformBufferArrayDynamicIndexing Bool32
	shaderSampledImageArrayDynamicIndexing  Bool32
	shaderStorageBufferArrayDynamicIndexing Bool32
	shaderStorageImageArrayDynamicIndexing  Bool32
	shaderClipDistance                      Bool32
	shaderCullDistance                      Bool32
	shaderFloat64                           Bool32
	shaderInt64                             Bool32
	shaderInt16                             Bool32
	shaderResourceResidency                 Bool32
	shaderResourceMinLod                    Bool32
	sparseBinding                           Bool32
	sparseResidencyBuffer                   Bool32
	sparseResidencyImage2D                  Bool32
	sparseResidencyImage3D                  Bool32
	sparseResidency2Samples                 Bool32
	sparseResidency4Samples                 Bool32
	sparseResidency8Samples                 Bool32
	sparseResidency16Samples                Bool32
	sparseResidencyAliased                  Bool32
	variableMultisampleRate                 Bool32
	inheritedQueries                        Bool32
}

pub type PhysicalDeviceLimits = C.VkPhysicalDeviceLimits

@[typedef]
pub struct C.VkPhysicalDeviceLimits {
pub mut:
	maxImageDimension1D                             u32
	maxImageDimension2D                             u32
	maxImageDimension3D                             u32
	maxImageDimensionCube                           u32
	maxImageArrayLayers                             u32
	maxTexelBufferElements                          u32
	maxUniformBufferRange                           u32
	maxStorageBufferRange                           u32
	maxPushConstantsSize                            u32
	maxMemoryAllocationCount                        u32
	maxSamplerAllocationCount                       u32
	bufferImageGranularity                          DeviceSize
	sparseAddressSpaceSize                          DeviceSize
	maxBoundDescriptorSets                          u32
	maxPerStageDescriptorSamplers                   u32
	maxPerStageDescriptorUniformBuffers             u32
	maxPerStageDescriptorStorageBuffers             u32
	maxPerStageDescriptorSampledImages              u32
	maxPerStageDescriptorStorageImages              u32
	maxPerStageDescriptorInputAttachments           u32
	maxPerStageResources                            u32
	maxDescriptorSetSamplers                        u32
	maxDescriptorSetUniformBuffers                  u32
	maxDescriptorSetUniformBuffersDynamic           u32
	maxDescriptorSetStorageBuffers                  u32
	maxDescriptorSetStorageBuffersDynamic           u32
	maxDescriptorSetSampledImages                   u32
	maxDescriptorSetStorageImages                   u32
	maxDescriptorSetInputAttachments                u32
	maxVertexInputAttributes                        u32
	maxVertexInputBindings                          u32
	maxVertexInputAttributeOffset                   u32
	maxVertexInputBindingStride                     u32
	maxVertexOutputComponents                       u32
	maxTessellationGenerationLevel                  u32
	maxTessellationPatchSize                        u32
	maxTessellationControlPerVertexInputComponents  u32
	maxTessellationControlPerVertexOutputComponents u32
	maxTessellationControlPerPatchOutputComponents  u32
	maxTessellationControlTotalOutputComponents     u32
	maxTessellationEvaluationInputComponents        u32
	maxTessellationEvaluationOutputComponents       u32
	maxGeometryShaderInvocations                    u32
	maxGeometryInputComponents                      u32
	maxGeometryOutputComponents                     u32
	maxGeometryOutputVertices                       u32
	maxGeometryTotalOutputComponents                u32
	maxFragmentInputComponents                      u32
	maxFragmentOutputAttachments                    u32
	maxFragmentDualSrcAttachments                   u32
	maxFragmentCombinedOutputResources              u32
	maxComputeSharedMemorySize                      u32
	maxComputeWorkGroupCount                        [3]u32
	maxComputeWorkGroupInvocations                  u32
	maxComputeWorkGroupSize                         [3]u32
	subPixelPrecisionBits                           u32
	subTexelPrecisionBits                           u32
	mipmapPrecisionBits                             u32
	maxDrawIndexedIndexValue                        u32
	maxDrawIndirectCount                            u32
	maxSamplerLodBias                               f32
	maxSamplerAnisotropy                            f32
	maxViewports                                    u32
	maxViewportDimensions                           [2]u32
	viewportBoundsRange                             [2]f32
	viewportSubPixelBits                            u32
	minMemoryMapAlignment                           usize
	minTexelBufferOffsetAlignment                   DeviceSize
	minUniformBufferOffsetAlignment                 DeviceSize
	minStorageBufferOffsetAlignment                 DeviceSize
	minTexelOffset                                  i32
	maxTexelOffset                                  u32
	minTexelGatherOffset                            i32
	maxTexelGatherOffset                            u32
	minInterpolationOffset                          f32
	maxInterpolationOffset                          f32
	subPixelInterpolationOffsetBits                 u32
	maxFramebufferWidth                             u32
	maxFramebufferHeight                            u32
	maxFramebufferLayers                            u32
	framebufferColorSampleCounts                    SampleCountFlags
	framebufferDepthSampleCounts                    SampleCountFlags
	framebufferStencilSampleCounts                  SampleCountFlags
	framebufferNoAttachmentsSampleCounts            SampleCountFlags
	maxColorAttachments                             u32
	sampledImageColorSampleCounts                   SampleCountFlags
	sampledImageIntegerSampleCounts                 SampleCountFlags
	sampledImageDepthSampleCounts                   SampleCountFlags
	sampledImageStencilSampleCounts                 SampleCountFlags
	storageImageSampleCounts                        SampleCountFlags
	maxSampleMaskWords                              u32
	timestampComputeAndGraphics                     Bool32
	timestampPeriod                                 f32
	maxClipDistances                                u32
	maxCullDistances                                u32
	maxCombinedClipAndCullDistances                 u32
	discreteQueuePriorities                         u32
	pointSizeRange                                  [2]f32
	lineWidthRange                                  [2]f32
	pointSizeGranularity                            f32
	lineWidthGranularity                            f32
	strictLines                                     Bool32
	standardSampleLocations                         Bool32
	optimalBufferCopyOffsetAlignment                DeviceSize
	optimalBufferCopyRowPitchAlignment              DeviceSize
	nonCoherentAtomSize                             DeviceSize
}

pub type PhysicalDeviceMemoryProperties = C.VkPhysicalDeviceMemoryProperties

@[typedef]
pub struct C.VkPhysicalDeviceMemoryProperties {
pub mut:
	memoryTypeCount u32
	memoryTypes     [max_memory_types]MemoryType
	memoryHeapCount u32
	memoryHeaps     [max_memory_heaps]MemoryHeap
}

pub type PhysicalDeviceSparseProperties = C.VkPhysicalDeviceSparseProperties

@[typedef]
pub struct C.VkPhysicalDeviceSparseProperties {
pub mut:
	residencyStandard2DBlockShape            Bool32
	residencyStandard2DMultisampleBlockShape Bool32
	residencyStandard3DBlockShape            Bool32
	residencyAlignedMipSize                  Bool32
	residencyNonResidentStrict               Bool32
}

pub type PhysicalDeviceProperties = C.VkPhysicalDeviceProperties

@[typedef]
pub struct C.VkPhysicalDeviceProperties {
pub mut:
	apiVersion        u32
	driverVersion     u32
	vendorID          u32
	deviceID          u32
	deviceType        PhysicalDeviceType
	deviceName        [max_physical_device_name_size]char
	pipelineCacheUUID [uuid_size]u8
	limits            PhysicalDeviceLimits
	sparseProperties  PhysicalDeviceSparseProperties
}

pub type QueueFamilyProperties = C.VkQueueFamilyProperties

@[typedef]
pub struct C.VkQueueFamilyProperties {
pub mut:
	queueFlags                  QueueFlags
	queueCount                  u32
	timestampValidBits          u32
	minImageTransferGranularity Extent3D
}

pub type DeviceQueueCreateInfo = C.VkDeviceQueueCreateInfo

@[typedef]
pub struct C.VkDeviceQueueCreateInfo {
pub mut:
	sType            StructureType = StructureType.device_queue_create_info
	pNext            voidptr       = unsafe { nil }
	flags            DeviceQueueCreateFlags
	queueFamilyIndex u32
	queueCount       u32
	pQueuePriorities &f32
}

pub type DeviceCreateInfo = C.VkDeviceCreateInfo

@[typedef]
pub struct C.VkDeviceCreateInfo {
pub mut:
	sType                StructureType = StructureType.device_create_info
	pNext                voidptr       = unsafe { nil }
	flags                DeviceCreateFlags
	queueCreateInfoCount u32
	pQueueCreateInfos    &DeviceQueueCreateInfo
	// enabledLayerCount is deprecated and should not be used
	enabledLayerCount u32
	// ppEnabledLayerNames is deprecated and should not be used
	ppEnabledLayerNames     &&char
	enabledExtensionCount   u32
	ppEnabledExtensionNames &&char
	pEnabledFeatures        &PhysicalDeviceFeatures
}

pub type ExtensionProperties = C.VkExtensionProperties

@[typedef]
pub struct C.VkExtensionProperties {
pub mut:
	extensionName [max_extension_name_size]char
	specVersion   u32
}

pub type LayerProperties = C.VkLayerProperties

@[typedef]
pub struct C.VkLayerProperties {
pub mut:
	layerName             [max_extension_name_size]char
	specVersion           u32
	implementationVersion u32
	description           [max_description_size]char
}

pub type SubmitInfo = C.VkSubmitInfo

@[typedef]
pub struct C.VkSubmitInfo {
pub mut:
	sType                StructureType = StructureType.submit_info
	pNext                voidptr       = unsafe { nil }
	waitSemaphoreCount   u32
	pWaitSemaphores      &Semaphore
	pWaitDstStageMask    &PipelineStageFlags
	commandBufferCount   u32
	pCommandBuffers      &CommandBuffer
	signalSemaphoreCount u32
	pSignalSemaphores    &Semaphore
}

pub type MappedMemoryRange = C.VkMappedMemoryRange

@[typedef]
pub struct C.VkMappedMemoryRange {
pub mut:
	sType  StructureType = StructureType.mapped_memory_range
	pNext  voidptr       = unsafe { nil }
	memory DeviceMemory
	offset DeviceSize
	size   DeviceSize
}

pub type MemoryAllocateInfo = C.VkMemoryAllocateInfo

@[typedef]
pub struct C.VkMemoryAllocateInfo {
pub mut:
	sType           StructureType = StructureType.memory_allocate_info
	pNext           voidptr       = unsafe { nil }
	allocationSize  DeviceSize
	memoryTypeIndex u32
}

pub type MemoryRequirements = C.VkMemoryRequirements

@[typedef]
pub struct C.VkMemoryRequirements {
pub mut:
	size           DeviceSize
	alignment      DeviceSize
	memoryTypeBits u32
}

pub type SparseMemoryBind = C.VkSparseMemoryBind

@[typedef]
pub struct C.VkSparseMemoryBind {
pub mut:
	resourceOffset DeviceSize
	size           DeviceSize
	memory         DeviceMemory
	memoryOffset   DeviceSize
	flags          SparseMemoryBindFlags
}

pub type SparseBufferMemoryBindInfo = C.VkSparseBufferMemoryBindInfo

@[typedef]
pub struct C.VkSparseBufferMemoryBindInfo {
pub mut:
	buffer    Buffer
	bindCount u32
	pBinds    &SparseMemoryBind
}

pub type SparseImageOpaqueMemoryBindInfo = C.VkSparseImageOpaqueMemoryBindInfo

@[typedef]
pub struct C.VkSparseImageOpaqueMemoryBindInfo {
pub mut:
	image     Image
	bindCount u32
	pBinds    &SparseMemoryBind
}

pub type ImageSubresource = C.VkImageSubresource

@[typedef]
pub struct C.VkImageSubresource {
pub mut:
	aspectMask ImageAspectFlags
	mipLevel   u32
	arrayLayer u32
}

pub type SparseImageMemoryBind = C.VkSparseImageMemoryBind

@[typedef]
pub struct C.VkSparseImageMemoryBind {
pub mut:
	subresource  ImageSubresource
	offset       Offset3D
	extent       Extent3D
	memory       DeviceMemory
	memoryOffset DeviceSize
	flags        SparseMemoryBindFlags
}

pub type SparseImageMemoryBindInfo = C.VkSparseImageMemoryBindInfo

@[typedef]
pub struct C.VkSparseImageMemoryBindInfo {
pub mut:
	image     Image
	bindCount u32
	pBinds    &SparseImageMemoryBind
}

pub type BindSparseInfo = C.VkBindSparseInfo

@[typedef]
pub struct C.VkBindSparseInfo {
pub mut:
	sType                StructureType = StructureType.bind_sparse_info
	pNext                voidptr       = unsafe { nil }
	waitSemaphoreCount   u32
	pWaitSemaphores      &Semaphore
	bufferBindCount      u32
	pBufferBinds         &SparseBufferMemoryBindInfo
	imageOpaqueBindCount u32
	pImageOpaqueBinds    &SparseImageOpaqueMemoryBindInfo
	imageBindCount       u32
	pImageBinds          &SparseImageMemoryBindInfo
	signalSemaphoreCount u32
	pSignalSemaphores    &Semaphore
}

pub type SparseImageFormatProperties = C.VkSparseImageFormatProperties

@[typedef]
pub struct C.VkSparseImageFormatProperties {
pub mut:
	aspectMask       ImageAspectFlags
	imageGranularity Extent3D
	flags            SparseImageFormatFlags
}

pub type SparseImageMemoryRequirements = C.VkSparseImageMemoryRequirements

@[typedef]
pub struct C.VkSparseImageMemoryRequirements {
pub mut:
	formatProperties     SparseImageFormatProperties
	imageMipTailFirstLod u32
	imageMipTailSize     DeviceSize
	imageMipTailOffset   DeviceSize
	imageMipTailStride   DeviceSize
}

pub type FenceCreateInfo = C.VkFenceCreateInfo

@[typedef]
pub struct C.VkFenceCreateInfo {
pub mut:
	sType StructureType = StructureType.fence_create_info
	pNext voidptr       = unsafe { nil }
	flags FenceCreateFlags
}

pub type SemaphoreCreateInfo = C.VkSemaphoreCreateInfo

@[typedef]
pub struct C.VkSemaphoreCreateInfo {
pub mut:
	sType StructureType = StructureType.semaphore_create_info
	pNext voidptr       = unsafe { nil }
	flags SemaphoreCreateFlags
}

pub type QueryPoolCreateInfo = C.VkQueryPoolCreateInfo

@[typedef]
pub struct C.VkQueryPoolCreateInfo {
pub mut:
	sType              StructureType = StructureType.query_pool_create_info
	pNext              voidptr       = unsafe { nil }
	flags              QueryPoolCreateFlags
	queryType          QueryType
	queryCount         u32
	pipelineStatistics QueryPipelineStatisticFlags
}

pub type BufferCreateInfo = C.VkBufferCreateInfo

@[typedef]
pub struct C.VkBufferCreateInfo {
pub mut:
	sType                 StructureType = StructureType.buffer_create_info
	pNext                 voidptr       = unsafe { nil }
	flags                 BufferCreateFlags
	size                  DeviceSize
	usage                 BufferUsageFlags
	sharingMode           SharingMode
	queueFamilyIndexCount u32
	pQueueFamilyIndices   &u32
}

pub type ImageCreateInfo = C.VkImageCreateInfo

@[typedef]
pub struct C.VkImageCreateInfo {
pub mut:
	sType                 StructureType = StructureType.image_create_info
	pNext                 voidptr       = unsafe { nil }
	flags                 ImageCreateFlags
	imageType             ImageType
	format                Format
	extent                Extent3D
	mipLevels             u32
	arrayLayers           u32
	samples               SampleCountFlagBits
	tiling                ImageTiling
	usage                 ImageUsageFlags
	sharingMode           SharingMode
	queueFamilyIndexCount u32
	pQueueFamilyIndices   &u32
	initialLayout         ImageLayout
}

pub type SubresourceLayout = C.VkSubresourceLayout

@[typedef]
pub struct C.VkSubresourceLayout {
pub mut:
	offset     DeviceSize
	size       DeviceSize
	rowPitch   DeviceSize
	arrayPitch DeviceSize
	depthPitch DeviceSize
}

pub type ComponentMapping = C.VkComponentMapping

@[typedef]
pub struct C.VkComponentMapping {
pub mut:
	r ComponentSwizzle
	g ComponentSwizzle
	b ComponentSwizzle
	a ComponentSwizzle
}

pub type ImageViewCreateInfo = C.VkImageViewCreateInfo

@[typedef]
pub struct C.VkImageViewCreateInfo {
pub mut:
	sType            StructureType = StructureType.image_view_create_info
	pNext            voidptr       = unsafe { nil }
	flags            ImageViewCreateFlags
	image            Image
	viewType         ImageViewType
	format           Format
	components       ComponentMapping
	subresourceRange ImageSubresourceRange
}

pub type CommandPoolCreateInfo = C.VkCommandPoolCreateInfo

@[typedef]
pub struct C.VkCommandPoolCreateInfo {
pub mut:
	sType            StructureType = StructureType.command_pool_create_info
	pNext            voidptr       = unsafe { nil }
	flags            CommandPoolCreateFlags
	queueFamilyIndex u32
}

pub type CommandBufferAllocateInfo = C.VkCommandBufferAllocateInfo

@[typedef]
pub struct C.VkCommandBufferAllocateInfo {
pub mut:
	sType              StructureType = StructureType.command_buffer_allocate_info
	pNext              voidptr       = unsafe { nil }
	commandPool        CommandPool
	level              CommandBufferLevel
	commandBufferCount u32
}

pub type CommandBufferInheritanceInfo = C.VkCommandBufferInheritanceInfo

@[typedef]
pub struct C.VkCommandBufferInheritanceInfo {
pub mut:
	sType                StructureType = StructureType.command_buffer_inheritance_info
	pNext                voidptr       = unsafe { nil }
	renderPass           RenderPass
	subpass              u32
	framebuffer          Framebuffer
	occlusionQueryEnable Bool32
	queryFlags           QueryControlFlags
	pipelineStatistics   QueryPipelineStatisticFlags
}

pub type CommandBufferBeginInfo = C.VkCommandBufferBeginInfo

@[typedef]
pub struct C.VkCommandBufferBeginInfo {
pub mut:
	sType            StructureType = StructureType.command_buffer_begin_info
	pNext            voidptr       = unsafe { nil }
	flags            CommandBufferUsageFlags
	pInheritanceInfo &CommandBufferInheritanceInfo
}

pub type BufferCopy = C.VkBufferCopy

@[typedef]
pub struct C.VkBufferCopy {
pub mut:
	srcOffset DeviceSize
	dstOffset DeviceSize
	size      DeviceSize
}

pub type ImageSubresourceLayers = C.VkImageSubresourceLayers

@[typedef]
pub struct C.VkImageSubresourceLayers {
pub mut:
	aspectMask     ImageAspectFlags
	mipLevel       u32
	baseArrayLayer u32
	layerCount     u32
}

pub type BufferImageCopy = C.VkBufferImageCopy

@[typedef]
pub struct C.VkBufferImageCopy {
pub mut:
	bufferOffset      DeviceSize
	bufferRowLength   u32
	bufferImageHeight u32
	imageSubresource  ImageSubresourceLayers
	imageOffset       Offset3D
	imageExtent       Extent3D
}

pub type ImageCopy = C.VkImageCopy

@[typedef]
pub struct C.VkImageCopy {
pub mut:
	srcSubresource ImageSubresourceLayers
	srcOffset      Offset3D
	dstSubresource ImageSubresourceLayers
	dstOffset      Offset3D
	extent         Extent3D
}

pub type DispatchIndirectCommand = C.VkDispatchIndirectCommand

@[typedef]
pub struct C.VkDispatchIndirectCommand {
pub mut:
	x u32
	y u32
	z u32
}

pub type PipelineCacheHeaderVersionOne = C.VkPipelineCacheHeaderVersionOne

@[typedef]
pub struct C.VkPipelineCacheHeaderVersionOne {
pub mut:
	headerSize        u32
	headerVersion     PipelineCacheHeaderVersion
	vendorID          u32
	deviceID          u32
	pipelineCacheUUID [uuid_size]u8
}

pub type EventCreateInfo = C.VkEventCreateInfo

@[typedef]
pub struct C.VkEventCreateInfo {
pub mut:
	sType StructureType = StructureType.event_create_info
	pNext voidptr       = unsafe { nil }
	flags EventCreateFlags
}

pub type BufferViewCreateInfo = C.VkBufferViewCreateInfo

@[typedef]
pub struct C.VkBufferViewCreateInfo {
pub mut:
	sType  StructureType = StructureType.buffer_view_create_info
	pNext  voidptr       = unsafe { nil }
	flags  BufferViewCreateFlags
	buffer Buffer
	format Format
	offset DeviceSize
	range  DeviceSize
}

// ShaderModuleCreateInfo extends VkPipelineShaderStageCreateInfo,VkDataGraphPipelineCreateInfoARM
pub type ShaderModuleCreateInfo = C.VkShaderModuleCreateInfo

@[typedef]
pub struct C.VkShaderModuleCreateInfo {
pub mut:
	sType    StructureType = StructureType.shader_module_create_info
	pNext    voidptr       = unsafe { nil }
	flags    ShaderModuleCreateFlags
	codeSize usize
	pCode    &u32
}

pub type PipelineCacheCreateInfo = C.VkPipelineCacheCreateInfo

@[typedef]
pub struct C.VkPipelineCacheCreateInfo {
pub mut:
	sType           StructureType = StructureType.pipeline_cache_create_info
	pNext           voidptr       = unsafe { nil }
	flags           PipelineCacheCreateFlags
	initialDataSize usize
	pInitialData    voidptr
}

pub type SpecializationMapEntry = C.VkSpecializationMapEntry

@[typedef]
pub struct C.VkSpecializationMapEntry {
pub mut:
	constantID u32
	offset     u32
	size       usize
}

pub type SpecializationInfo = C.VkSpecializationInfo

@[typedef]
pub struct C.VkSpecializationInfo {
pub mut:
	mapEntryCount u32
	pMapEntries   &SpecializationMapEntry
	dataSize      usize
	pData         voidptr
}

pub type PipelineShaderStageCreateInfo = C.VkPipelineShaderStageCreateInfo

@[typedef]
pub struct C.VkPipelineShaderStageCreateInfo {
pub mut:
	sType               StructureType = StructureType.pipeline_shader_stage_create_info
	pNext               voidptr       = unsafe { nil }
	flags               PipelineShaderStageCreateFlags
	stage               ShaderStageFlagBits
	module              ShaderModule
	pName               &char
	pSpecializationInfo &SpecializationInfo
}

pub type ComputePipelineCreateInfo = C.VkComputePipelineCreateInfo

@[typedef]
pub struct C.VkComputePipelineCreateInfo {
pub mut:
	sType              StructureType = StructureType.compute_pipeline_create_info
	pNext              voidptr       = unsafe { nil }
	flags              PipelineCreateFlags
	stage              PipelineShaderStageCreateInfo
	layout             PipelineLayout
	basePipelineHandle Pipeline
	basePipelineIndex  i32
}

pub type PushConstantRange = C.VkPushConstantRange

@[typedef]
pub struct C.VkPushConstantRange {
pub mut:
	stageFlags ShaderStageFlags
	offset     u32
	size       u32
}

// PipelineLayoutCreateInfo extends VkBindDescriptorSetsInfo,VkPushConstantsInfo,VkPushDescriptorSetInfo,VkPushDescriptorSetWithTemplateInfo,VkSetDescriptorBufferOffsetsInfoEXT,VkBindDescriptorBufferEmbeddedSamplersInfoEXT,VkIndirectCommandsLayoutCreateInfoEXT
pub type PipelineLayoutCreateInfo = C.VkPipelineLayoutCreateInfo

@[typedef]
pub struct C.VkPipelineLayoutCreateInfo {
pub mut:
	sType                  StructureType = StructureType.pipeline_layout_create_info
	pNext                  voidptr       = unsafe { nil }
	flags                  PipelineLayoutCreateFlags
	setLayoutCount         u32
	pSetLayouts            &DescriptorSetLayout
	pushConstantRangeCount u32
	pPushConstantRanges    &PushConstantRange
}

pub type SamplerCreateInfo = C.VkSamplerCreateInfo

@[typedef]
pub struct C.VkSamplerCreateInfo {
pub mut:
	sType                   StructureType = StructureType.sampler_create_info
	pNext                   voidptr       = unsafe { nil }
	flags                   SamplerCreateFlags
	magFilter               Filter
	minFilter               Filter
	mipmapMode              SamplerMipmapMode
	addressModeU            SamplerAddressMode
	addressModeV            SamplerAddressMode
	addressModeW            SamplerAddressMode
	mipLodBias              f32
	anisotropyEnable        Bool32
	maxAnisotropy           f32
	compareEnable           Bool32
	compareOp               CompareOp
	minLod                  f32
	maxLod                  f32
	borderColor             BorderColor
	unnormalizedCoordinates Bool32
}

pub type CopyDescriptorSet = C.VkCopyDescriptorSet

@[typedef]
pub struct C.VkCopyDescriptorSet {
pub mut:
	sType           StructureType = StructureType.copy_descriptor_set
	pNext           voidptr       = unsafe { nil }
	srcSet          DescriptorSet
	srcBinding      u32
	srcArrayElement u32
	dstSet          DescriptorSet
	dstBinding      u32
	dstArrayElement u32
	descriptorCount u32
}

pub type DescriptorBufferInfo = C.VkDescriptorBufferInfo

@[typedef]
pub struct C.VkDescriptorBufferInfo {
pub mut:
	buffer Buffer
	offset DeviceSize
	range  DeviceSize
}

pub type DescriptorImageInfo = C.VkDescriptorImageInfo

@[typedef]
pub struct C.VkDescriptorImageInfo {
pub mut:
	sampler     Sampler
	imageView   ImageView
	imageLayout ImageLayout
}

pub type DescriptorPoolSize = C.VkDescriptorPoolSize

@[typedef]
pub struct C.VkDescriptorPoolSize {
pub mut:
	type            DescriptorType
	descriptorCount u32
}

pub type DescriptorPoolCreateInfo = C.VkDescriptorPoolCreateInfo

@[typedef]
pub struct C.VkDescriptorPoolCreateInfo {
pub mut:
	sType         StructureType = StructureType.descriptor_pool_create_info
	pNext         voidptr       = unsafe { nil }
	flags         DescriptorPoolCreateFlags
	maxSets       u32
	poolSizeCount u32
	pPoolSizes    &DescriptorPoolSize
}

pub type DescriptorSetAllocateInfo = C.VkDescriptorSetAllocateInfo

@[typedef]
pub struct C.VkDescriptorSetAllocateInfo {
pub mut:
	sType              StructureType = StructureType.descriptor_set_allocate_info
	pNext              voidptr       = unsafe { nil }
	descriptorPool     DescriptorPool
	descriptorSetCount u32
	pSetLayouts        &DescriptorSetLayout
}

pub type DescriptorSetLayoutBinding = C.VkDescriptorSetLayoutBinding

@[typedef]
pub struct C.VkDescriptorSetLayoutBinding {
pub mut:
	binding            u32
	descriptorType     DescriptorType
	descriptorCount    u32
	stageFlags         ShaderStageFlags
	pImmutableSamplers &Sampler
}

pub type DescriptorSetLayoutCreateInfo = C.VkDescriptorSetLayoutCreateInfo

@[typedef]
pub struct C.VkDescriptorSetLayoutCreateInfo {
pub mut:
	sType        StructureType = StructureType.descriptor_set_layout_create_info
	pNext        voidptr       = unsafe { nil }
	flags        DescriptorSetLayoutCreateFlags
	bindingCount u32
	pBindings    &DescriptorSetLayoutBinding
}

pub type WriteDescriptorSet = C.VkWriteDescriptorSet

@[typedef]
pub struct C.VkWriteDescriptorSet {
pub mut:
	sType            StructureType = StructureType.write_descriptor_set
	pNext            voidptr       = unsafe { nil }
	dstSet           DescriptorSet
	dstBinding       u32
	dstArrayElement  u32
	descriptorCount  u32
	descriptorType   DescriptorType
	pImageInfo       &DescriptorImageInfo
	pBufferInfo      &DescriptorBufferInfo
	pTexelBufferView &BufferView
}

pub type ClearColorValue = C.VkClearColorValue

@[typedef]
pub union C.VkClearColorValue {
pub mut:
	float32 [4]f32
	int32   [4]i32
	uint32  [4]u32
}

pub type DrawIndexedIndirectCommand = C.VkDrawIndexedIndirectCommand

@[typedef]
pub struct C.VkDrawIndexedIndirectCommand {
pub mut:
	indexCount    u32
	instanceCount u32
	firstIndex    u32
	vertexOffset  i32
	firstInstance u32
}

pub type DrawIndirectCommand = C.VkDrawIndirectCommand

@[typedef]
pub struct C.VkDrawIndirectCommand {
pub mut:
	vertexCount   u32
	instanceCount u32
	firstVertex   u32
	firstInstance u32
}

pub type VertexInputBindingDescription = C.VkVertexInputBindingDescription

@[typedef]
pub struct C.VkVertexInputBindingDescription {
pub mut:
	binding   u32
	stride    u32
	inputRate VertexInputRate
}

pub type VertexInputAttributeDescription = C.VkVertexInputAttributeDescription

@[typedef]
pub struct C.VkVertexInputAttributeDescription {
pub mut:
	location u32
	binding  u32
	format   Format
	offset   u32
}

pub type PipelineVertexInputStateCreateInfo = C.VkPipelineVertexInputStateCreateInfo

@[typedef]
pub struct C.VkPipelineVertexInputStateCreateInfo {
pub mut:
	sType                           StructureType = StructureType.pipeline_vertex_input_state_create_info
	pNext                           voidptr       = unsafe { nil }
	flags                           PipelineVertexInputStateCreateFlags
	vertexBindingDescriptionCount   u32
	pVertexBindingDescriptions      &VertexInputBindingDescription
	vertexAttributeDescriptionCount u32
	pVertexAttributeDescriptions    &VertexInputAttributeDescription
}

pub type PipelineInputAssemblyStateCreateInfo = C.VkPipelineInputAssemblyStateCreateInfo

@[typedef]
pub struct C.VkPipelineInputAssemblyStateCreateInfo {
pub mut:
	sType                  StructureType = StructureType.pipeline_input_assembly_state_create_info
	pNext                  voidptr       = unsafe { nil }
	flags                  PipelineInputAssemblyStateCreateFlags
	topology               PrimitiveTopology
	primitiveRestartEnable Bool32
}

pub type PipelineTessellationStateCreateInfo = C.VkPipelineTessellationStateCreateInfo

@[typedef]
pub struct C.VkPipelineTessellationStateCreateInfo {
pub mut:
	sType              StructureType = StructureType.pipeline_tessellation_state_create_info
	pNext              voidptr       = unsafe { nil }
	flags              PipelineTessellationStateCreateFlags
	patchControlPoints u32
}

pub type Viewport = C.VkViewport

@[typedef]
pub struct C.VkViewport {
pub mut:
	x        f32
	y        f32
	width    f32
	height   f32
	minDepth f32
	maxDepth f32
}

pub type PipelineViewportStateCreateInfo = C.VkPipelineViewportStateCreateInfo

@[typedef]
pub struct C.VkPipelineViewportStateCreateInfo {
pub mut:
	sType         StructureType = StructureType.pipeline_viewport_state_create_info
	pNext         voidptr       = unsafe { nil }
	flags         PipelineViewportStateCreateFlags
	viewportCount u32
	pViewports    &Viewport
	scissorCount  u32
	pScissors     &Rect2D
}

pub type PipelineRasterizationStateCreateInfo = C.VkPipelineRasterizationStateCreateInfo

@[typedef]
pub struct C.VkPipelineRasterizationStateCreateInfo {
pub mut:
	sType                   StructureType = StructureType.pipeline_rasterization_state_create_info
	pNext                   voidptr       = unsafe { nil }
	flags                   PipelineRasterizationStateCreateFlags
	depthClampEnable        Bool32
	rasterizerDiscardEnable Bool32
	polygonMode             PolygonMode
	cullMode                CullModeFlags
	frontFace               FrontFace
	depthBiasEnable         Bool32
	depthBiasConstantFactor f32
	depthBiasClamp          f32
	depthBiasSlopeFactor    f32
	lineWidth               f32
}

pub type PipelineMultisampleStateCreateInfo = C.VkPipelineMultisampleStateCreateInfo

@[typedef]
pub struct C.VkPipelineMultisampleStateCreateInfo {
pub mut:
	sType                 StructureType = StructureType.pipeline_multisample_state_create_info
	pNext                 voidptr       = unsafe { nil }
	flags                 PipelineMultisampleStateCreateFlags
	rasterizationSamples  SampleCountFlagBits
	sampleShadingEnable   Bool32
	minSampleShading      f32
	pSampleMask           &SampleMask
	alphaToCoverageEnable Bool32
	alphaToOneEnable      Bool32
}

pub type StencilOpState = C.VkStencilOpState

@[typedef]
pub struct C.VkStencilOpState {
pub mut:
	failOp      StencilOp
	passOp      StencilOp
	depthFailOp StencilOp
	compareOp   CompareOp
	compareMask u32
	writeMask   u32
	reference   u32
}

pub type PipelineDepthStencilStateCreateInfo = C.VkPipelineDepthStencilStateCreateInfo

@[typedef]
pub struct C.VkPipelineDepthStencilStateCreateInfo {
pub mut:
	sType                 StructureType = StructureType.pipeline_depth_stencil_state_create_info
	pNext                 voidptr       = unsafe { nil }
	flags                 PipelineDepthStencilStateCreateFlags
	depthTestEnable       Bool32
	depthWriteEnable      Bool32
	depthCompareOp        CompareOp
	depthBoundsTestEnable Bool32
	stencilTestEnable     Bool32
	front                 StencilOpState
	back                  StencilOpState
	minDepthBounds        f32
	maxDepthBounds        f32
}

pub type PipelineColorBlendAttachmentState = C.VkPipelineColorBlendAttachmentState

@[typedef]
pub struct C.VkPipelineColorBlendAttachmentState {
pub mut:
	blendEnable         Bool32
	srcColorBlendFactor BlendFactor
	dstColorBlendFactor BlendFactor
	colorBlendOp        BlendOp
	srcAlphaBlendFactor BlendFactor
	dstAlphaBlendFactor BlendFactor
	alphaBlendOp        BlendOp
	colorWriteMask      ColorComponentFlags
}

pub type PipelineColorBlendStateCreateInfo = C.VkPipelineColorBlendStateCreateInfo

@[typedef]
pub struct C.VkPipelineColorBlendStateCreateInfo {
pub mut:
	sType           StructureType = StructureType.pipeline_color_blend_state_create_info
	pNext           voidptr       = unsafe { nil }
	flags           PipelineColorBlendStateCreateFlags
	logicOpEnable   Bool32
	logicOp         LogicOp
	attachmentCount u32
	pAttachments    &PipelineColorBlendAttachmentState
	blendConstants  [4]f32
}

pub type PipelineDynamicStateCreateInfo = C.VkPipelineDynamicStateCreateInfo

@[typedef]
pub struct C.VkPipelineDynamicStateCreateInfo {
pub mut:
	sType             StructureType = StructureType.pipeline_dynamic_state_create_info
	pNext             voidptr       = unsafe { nil }
	flags             PipelineDynamicStateCreateFlags
	dynamicStateCount u32
	pDynamicStates    &DynamicState
}

pub type GraphicsPipelineCreateInfo = C.VkGraphicsPipelineCreateInfo

@[typedef]
pub struct C.VkGraphicsPipelineCreateInfo {
pub mut:
	sType               StructureType = StructureType.graphics_pipeline_create_info
	pNext               voidptr       = unsafe { nil }
	flags               PipelineCreateFlags
	stageCount          u32
	pStages             &PipelineShaderStageCreateInfo
	pVertexInputState   &PipelineVertexInputStateCreateInfo
	pInputAssemblyState &PipelineInputAssemblyStateCreateInfo
	pTessellationState  &PipelineTessellationStateCreateInfo
	pViewportState      &PipelineViewportStateCreateInfo
	pRasterizationState &PipelineRasterizationStateCreateInfo
	pMultisampleState   &PipelineMultisampleStateCreateInfo
	pDepthStencilState  &PipelineDepthStencilStateCreateInfo
	pColorBlendState    &PipelineColorBlendStateCreateInfo
	pDynamicState       &PipelineDynamicStateCreateInfo
	layout              PipelineLayout
	renderPass          RenderPass
	subpass             u32
	basePipelineHandle  Pipeline
	basePipelineIndex   i32
}

pub type AttachmentDescription = C.VkAttachmentDescription

@[typedef]
pub struct C.VkAttachmentDescription {
pub mut:
	flags          AttachmentDescriptionFlags
	format         Format
	samples        SampleCountFlagBits
	loadOp         AttachmentLoadOp
	storeOp        AttachmentStoreOp
	stencilLoadOp  AttachmentLoadOp
	stencilStoreOp AttachmentStoreOp
	initialLayout  ImageLayout
	finalLayout    ImageLayout
}

pub type AttachmentReference = C.VkAttachmentReference

@[typedef]
pub struct C.VkAttachmentReference {
pub mut:
	attachment u32
	layout     ImageLayout
}

pub type FramebufferCreateInfo = C.VkFramebufferCreateInfo

@[typedef]
pub struct C.VkFramebufferCreateInfo {
pub mut:
	sType           StructureType = StructureType.framebuffer_create_info
	pNext           voidptr       = unsafe { nil }
	flags           FramebufferCreateFlags
	renderPass      RenderPass
	attachmentCount u32
	pAttachments    &ImageView
	width           u32
	height          u32
	layers          u32
}

pub type SubpassDescription = C.VkSubpassDescription

@[typedef]
pub struct C.VkSubpassDescription {
pub mut:
	flags                   SubpassDescriptionFlags
	pipelineBindPoint       PipelineBindPoint
	inputAttachmentCount    u32
	pInputAttachments       &AttachmentReference
	colorAttachmentCount    u32
	pColorAttachments       &AttachmentReference
	pResolveAttachments     &AttachmentReference
	pDepthStencilAttachment &AttachmentReference
	preserveAttachmentCount u32
	pPreserveAttachments    &u32
}

pub type SubpassDependency = C.VkSubpassDependency

@[typedef]
pub struct C.VkSubpassDependency {
pub mut:
	srcSubpass      u32
	dstSubpass      u32
	srcStageMask    PipelineStageFlags
	dstStageMask    PipelineStageFlags
	srcAccessMask   AccessFlags
	dstAccessMask   AccessFlags
	dependencyFlags DependencyFlags
}

pub type RenderPassCreateInfo = C.VkRenderPassCreateInfo

@[typedef]
pub struct C.VkRenderPassCreateInfo {
pub mut:
	sType           StructureType = StructureType.render_pass_create_info
	pNext           voidptr       = unsafe { nil }
	flags           RenderPassCreateFlags
	attachmentCount u32
	pAttachments    &AttachmentDescription
	subpassCount    u32
	pSubpasses      &SubpassDescription
	dependencyCount u32
	pDependencies   &SubpassDependency
}

pub type ClearDepthStencilValue = C.VkClearDepthStencilValue

@[typedef]
pub struct C.VkClearDepthStencilValue {
pub mut:
	depth   f32
	stencil u32
}

pub type ClearValue = C.VkClearValue

@[typedef]
pub union C.VkClearValue {
pub mut:
	color        ClearColorValue
	depthStencil ClearDepthStencilValue
}

pub type ClearAttachment = C.VkClearAttachment

@[typedef]
pub struct C.VkClearAttachment {
pub mut:
	aspectMask      ImageAspectFlags
	colorAttachment u32
	clearValue      ClearValue
}

pub type ClearRect = C.VkClearRect

@[typedef]
pub struct C.VkClearRect {
pub mut:
	rect           Rect2D
	baseArrayLayer u32
	layerCount     u32
}

pub type ImageBlit = C.VkImageBlit

@[typedef]
pub struct C.VkImageBlit {
pub mut:
	srcSubresource ImageSubresourceLayers
	srcOffsets     [2]Offset3D
	dstSubresource ImageSubresourceLayers
	dstOffsets     [2]Offset3D
}

pub type ImageResolve = C.VkImageResolve

@[typedef]
pub struct C.VkImageResolve {
pub mut:
	srcSubresource ImageSubresourceLayers
	srcOffset      Offset3D
	dstSubresource ImageSubresourceLayers
	dstOffset      Offset3D
	extent         Extent3D
}

pub type RenderPassBeginInfo = C.VkRenderPassBeginInfo

@[typedef]
pub struct C.VkRenderPassBeginInfo {
pub mut:
	sType           StructureType = StructureType.render_pass_begin_info
	pNext           voidptr       = unsafe { nil }
	renderPass      RenderPass
	framebuffer     Framebuffer
	renderArea      Rect2D
	clearValueCount u32
	pClearValues    &ClearValue
}

@[keep_args_alive]
fn C.vkCreateInstance(p_create_info &InstanceCreateInfo, p_allocator &AllocationCallbacks, p_instance &Instance) Result

pub type PFN_vkCreateInstance = fn (p_create_info &InstanceCreateInfo, p_allocator &AllocationCallbacks, p_instance &Instance) Result

@[inline]
pub fn create_instance(p_create_info &InstanceCreateInfo,
	p_allocator &AllocationCallbacks,
	p_instance &Instance) Result {
	return C.vkCreateInstance(p_create_info, p_allocator, p_instance)
}

@[keep_args_alive]
fn C.vkDestroyInstance(instance Instance, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyInstance = fn (instance Instance, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_instance(instance Instance,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyInstance(instance, p_allocator)
}

@[keep_args_alive]
fn C.vkEnumeratePhysicalDevices(instance Instance, p_physical_device_count &u32, p_physical_devices &PhysicalDevice) Result

pub type PFN_vkEnumeratePhysicalDevices = fn (instance Instance, p_physical_device_count &u32, p_physical_devices &PhysicalDevice) Result

@[inline]
pub fn enumerate_physical_devices(instance Instance,
	p_physical_device_count &u32,
	p_physical_devices &PhysicalDevice) Result {
	return C.vkEnumeratePhysicalDevices(instance, p_physical_device_count, p_physical_devices)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceFeatures(physical_device PhysicalDevice, mut p_features PhysicalDeviceFeatures)

pub type PFN_vkGetPhysicalDeviceFeatures = fn (physical_device PhysicalDevice, mut p_features PhysicalDeviceFeatures)

@[inline]
pub fn get_physical_device_features(physical_device PhysicalDevice,
	mut p_features PhysicalDeviceFeatures) {
	C.vkGetPhysicalDeviceFeatures(physical_device, mut p_features)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceFormatProperties(physical_device PhysicalDevice, format Format, mut p_format_properties FormatProperties)

pub type PFN_vkGetPhysicalDeviceFormatProperties = fn (physical_device PhysicalDevice, format Format, mut p_format_properties FormatProperties)

@[inline]
pub fn get_physical_device_format_properties(physical_device PhysicalDevice,
	format Format,
	mut p_format_properties FormatProperties) {
	C.vkGetPhysicalDeviceFormatProperties(physical_device, format, mut p_format_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceImageFormatProperties(physical_device PhysicalDevice, format Format, type_param ImageType, tiling ImageTiling, usage ImageUsageFlags, flags ImageCreateFlags, mut p_image_format_properties ImageFormatProperties) Result

pub type PFN_vkGetPhysicalDeviceImageFormatProperties = fn (physical_device PhysicalDevice, format Format, type_param ImageType, tiling ImageTiling, usage ImageUsageFlags, flags ImageCreateFlags, mut p_image_format_properties ImageFormatProperties) Result

@[inline]
pub fn get_physical_device_image_format_properties(physical_device PhysicalDevice,
	format Format,
	type_param ImageType,
	tiling ImageTiling,
	usage ImageUsageFlags,
	flags ImageCreateFlags,
	mut p_image_format_properties ImageFormatProperties) Result {
	return C.vkGetPhysicalDeviceImageFormatProperties(physical_device, format, type_param,
		tiling, usage, flags, mut p_image_format_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceProperties(physical_device PhysicalDevice, mut p_properties PhysicalDeviceProperties)

pub type PFN_vkGetPhysicalDeviceProperties = fn (physical_device PhysicalDevice, mut p_properties PhysicalDeviceProperties)

@[inline]
pub fn get_physical_device_properties(physical_device PhysicalDevice,
	mut p_properties PhysicalDeviceProperties) {
	C.vkGetPhysicalDeviceProperties(physical_device, mut p_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceQueueFamilyProperties(physical_device PhysicalDevice, p_queue_family_property_count &u32, mut p_queue_family_properties QueueFamilyProperties)

pub type PFN_vkGetPhysicalDeviceQueueFamilyProperties = fn (physical_device PhysicalDevice, p_queue_family_property_count &u32, mut p_queue_family_properties QueueFamilyProperties)

@[inline]
pub fn get_physical_device_queue_family_properties(physical_device PhysicalDevice,
	p_queue_family_property_count &u32,
	mut p_queue_family_properties QueueFamilyProperties) {
	C.vkGetPhysicalDeviceQueueFamilyProperties(physical_device, p_queue_family_property_count, mut
		p_queue_family_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceMemoryProperties(physical_device PhysicalDevice, mut p_memory_properties PhysicalDeviceMemoryProperties)

pub type PFN_vkGetPhysicalDeviceMemoryProperties = fn (physical_device PhysicalDevice, mut p_memory_properties PhysicalDeviceMemoryProperties)

@[inline]
pub fn get_physical_device_memory_properties(physical_device PhysicalDevice,
	mut p_memory_properties PhysicalDeviceMemoryProperties) {
	C.vkGetPhysicalDeviceMemoryProperties(physical_device, mut p_memory_properties)
}

@[keep_args_alive]
fn C.vkGetInstanceProcAddr(instance Instance, p_name &char) voidptr

pub type PFN_vkGetInstanceProcAddr = fn (instance Instance, p_name &char)

@[inline]
pub fn get_instance_proc_addr(instance Instance,
	p_name &char) voidptr {
	return C.vkGetInstanceProcAddr(instance, p_name)
}

@[keep_args_alive]
fn C.vkGetDeviceProcAddr(device Device, p_name &char) voidptr

pub type PFN_vkGetDeviceProcAddr = fn (device Device, p_name &char)

@[inline]
pub fn get_device_proc_addr(device Device,
	p_name &char) voidptr {
	return C.vkGetDeviceProcAddr(device, p_name)
}

@[keep_args_alive]
fn C.vkCreateDevice(physical_device PhysicalDevice, p_create_info &DeviceCreateInfo, p_allocator &AllocationCallbacks, p_device &Device) Result

pub type PFN_vkCreateDevice = fn (physical_device PhysicalDevice, p_create_info &DeviceCreateInfo, p_allocator &AllocationCallbacks, p_device &Device) Result

@[inline]
pub fn create_device(physical_device PhysicalDevice,
	p_create_info &DeviceCreateInfo,
	p_allocator &AllocationCallbacks,
	p_device &Device) Result {
	return C.vkCreateDevice(physical_device, p_create_info, p_allocator, p_device)
}

@[keep_args_alive]
fn C.vkDestroyDevice(device Device, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyDevice = fn (device Device, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_device(device Device,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyDevice(device, p_allocator)
}

@[keep_args_alive]
fn C.vkEnumerateInstanceExtensionProperties(p_layer_name &char, p_property_count &u32, mut p_properties ExtensionProperties) Result

pub type PFN_vkEnumerateInstanceExtensionProperties = fn (p_layer_name &char, p_property_count &u32, mut p_properties ExtensionProperties) Result

@[inline]
pub fn enumerate_instance_extension_properties(p_layer_name &char,
	p_property_count &u32,
	mut p_properties ExtensionProperties) Result {
	return C.vkEnumerateInstanceExtensionProperties(p_layer_name, p_property_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkEnumerateDeviceExtensionProperties(physical_device PhysicalDevice, p_layer_name &char, p_property_count &u32, mut p_properties ExtensionProperties) Result

pub type PFN_vkEnumerateDeviceExtensionProperties = fn (physical_device PhysicalDevice, p_layer_name &char, p_property_count &u32, mut p_properties ExtensionProperties) Result

@[inline]
pub fn enumerate_device_extension_properties(physical_device PhysicalDevice,
	p_layer_name &char,
	p_property_count &u32,
	mut p_properties ExtensionProperties) Result {
	return C.vkEnumerateDeviceExtensionProperties(physical_device, p_layer_name, p_property_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkEnumerateInstanceLayerProperties(p_property_count &u32, mut p_properties LayerProperties) Result

pub type PFN_vkEnumerateInstanceLayerProperties = fn (p_property_count &u32, mut p_properties LayerProperties) Result

@[inline]
pub fn enumerate_instance_layer_properties(p_property_count &u32,
	mut p_properties LayerProperties) Result {
	return C.vkEnumerateInstanceLayerProperties(p_property_count, mut p_properties)
}

@[keep_args_alive]
fn C.vkEnumerateDeviceLayerProperties(physical_device PhysicalDevice, p_property_count &u32, mut p_properties LayerProperties) Result

pub type PFN_vkEnumerateDeviceLayerProperties = fn (physical_device PhysicalDevice, p_property_count &u32, mut p_properties LayerProperties) Result

@[inline]
pub fn enumerate_device_layer_properties(physical_device PhysicalDevice,
	p_property_count &u32,
	mut p_properties LayerProperties) Result {
	return C.vkEnumerateDeviceLayerProperties(physical_device, p_property_count, mut p_properties)
}

@[keep_args_alive]
fn C.vkGetDeviceQueue(device Device, queue_family_index u32, queue_index u32, p_queue &Queue)

pub type PFN_vkGetDeviceQueue = fn (device Device, queue_family_index u32, queue_index u32, p_queue &Queue)

@[inline]
pub fn get_device_queue(device Device,
	queue_family_index u32,
	queue_index u32,
	p_queue &Queue) {
	C.vkGetDeviceQueue(device, queue_family_index, queue_index, p_queue)
}

@[keep_args_alive]
fn C.vkQueueSubmit(queue Queue, submit_count u32, p_submits &SubmitInfo, fence Fence) Result

pub type PFN_vkQueueSubmit = fn (queue Queue, submit_count u32, p_submits &SubmitInfo, fence Fence) Result

@[inline]
pub fn queue_submit(queue Queue,
	submit_count u32,
	p_submits &SubmitInfo,
	fence Fence) Result {
	return C.vkQueueSubmit(queue, submit_count, p_submits, fence)
}

@[keep_args_alive]
fn C.vkQueueWaitIdle(queue Queue) Result

pub type PFN_vkQueueWaitIdle = fn (queue Queue) Result

@[inline]
pub fn queue_wait_idle(queue Queue) Result {
	return C.vkQueueWaitIdle(queue)
}

@[keep_args_alive]
fn C.vkDeviceWaitIdle(device Device) Result

pub type PFN_vkDeviceWaitIdle = fn (device Device) Result

@[inline]
pub fn device_wait_idle(device Device) Result {
	return C.vkDeviceWaitIdle(device)
}

@[keep_args_alive]
fn C.vkAllocateMemory(device Device, p_allocate_info &MemoryAllocateInfo, p_allocator &AllocationCallbacks, p_memory &DeviceMemory) Result

pub type PFN_vkAllocateMemory = fn (device Device, p_allocate_info &MemoryAllocateInfo, p_allocator &AllocationCallbacks, p_memory &DeviceMemory) Result

@[inline]
pub fn allocate_memory(device Device,
	p_allocate_info &MemoryAllocateInfo,
	p_allocator &AllocationCallbacks,
	p_memory &DeviceMemory) Result {
	return C.vkAllocateMemory(device, p_allocate_info, p_allocator, p_memory)
}

@[keep_args_alive]
fn C.vkFreeMemory(device Device, memory DeviceMemory, p_allocator &AllocationCallbacks)

pub type PFN_vkFreeMemory = fn (device Device, memory DeviceMemory, p_allocator &AllocationCallbacks)

@[inline]
pub fn free_memory(device Device,
	memory DeviceMemory,
	p_allocator &AllocationCallbacks) {
	C.vkFreeMemory(device, memory, p_allocator)
}

@[keep_args_alive]
fn C.vkMapMemory(device Device, memory DeviceMemory, offset DeviceSize, size DeviceSize, flags MemoryMapFlags, pp_data &voidptr) Result

pub type PFN_vkMapMemory = fn (device Device, memory DeviceMemory, offset DeviceSize, size DeviceSize, flags MemoryMapFlags, pp_data &voidptr) Result

@[inline]
pub fn map_memory(device Device,
	memory DeviceMemory,
	offset DeviceSize,
	size DeviceSize,
	flags MemoryMapFlags,
	pp_data &voidptr) Result {
	return C.vkMapMemory(device, memory, offset, size, flags, pp_data)
}

@[keep_args_alive]
fn C.vkUnmapMemory(device Device, memory DeviceMemory)

pub type PFN_vkUnmapMemory = fn (device Device, memory DeviceMemory)

@[inline]
pub fn unmap_memory(device Device,
	memory DeviceMemory) {
	C.vkUnmapMemory(device, memory)
}

@[keep_args_alive]
fn C.vkFlushMappedMemoryRanges(device Device, memory_range_count u32, p_memory_ranges &MappedMemoryRange) Result

pub type PFN_vkFlushMappedMemoryRanges = fn (device Device, memory_range_count u32, p_memory_ranges &MappedMemoryRange) Result

@[inline]
pub fn flush_mapped_memory_ranges(device Device,
	memory_range_count u32,
	p_memory_ranges &MappedMemoryRange) Result {
	return C.vkFlushMappedMemoryRanges(device, memory_range_count, p_memory_ranges)
}

@[keep_args_alive]
fn C.vkInvalidateMappedMemoryRanges(device Device, memory_range_count u32, p_memory_ranges &MappedMemoryRange) Result

pub type PFN_vkInvalidateMappedMemoryRanges = fn (device Device, memory_range_count u32, p_memory_ranges &MappedMemoryRange) Result

@[inline]
pub fn invalidate_mapped_memory_ranges(device Device,
	memory_range_count u32,
	p_memory_ranges &MappedMemoryRange) Result {
	return C.vkInvalidateMappedMemoryRanges(device, memory_range_count, p_memory_ranges)
}

@[keep_args_alive]
fn C.vkGetDeviceMemoryCommitment(device Device, memory DeviceMemory, p_committed_memory_in_bytes &DeviceSize)

pub type PFN_vkGetDeviceMemoryCommitment = fn (device Device, memory DeviceMemory, p_committed_memory_in_bytes &DeviceSize)

@[inline]
pub fn get_device_memory_commitment(device Device,
	memory DeviceMemory,
	p_committed_memory_in_bytes &DeviceSize) {
	C.vkGetDeviceMemoryCommitment(device, memory, p_committed_memory_in_bytes)
}

@[keep_args_alive]
fn C.vkBindBufferMemory(device Device, buffer Buffer, memory DeviceMemory, memory_offset DeviceSize) Result

pub type PFN_vkBindBufferMemory = fn (device Device, buffer Buffer, memory DeviceMemory, memory_offset DeviceSize) Result

@[inline]
pub fn bind_buffer_memory(device Device,
	buffer Buffer,
	memory DeviceMemory,
	memory_offset DeviceSize) Result {
	return C.vkBindBufferMemory(device, buffer, memory, memory_offset)
}

@[keep_args_alive]
fn C.vkBindImageMemory(device Device, image Image, memory DeviceMemory, memory_offset DeviceSize) Result

pub type PFN_vkBindImageMemory = fn (device Device, image Image, memory DeviceMemory, memory_offset DeviceSize) Result

@[inline]
pub fn bind_image_memory(device Device,
	image Image,
	memory DeviceMemory,
	memory_offset DeviceSize) Result {
	return C.vkBindImageMemory(device, image, memory, memory_offset)
}

@[keep_args_alive]
fn C.vkGetBufferMemoryRequirements(device Device, buffer Buffer, mut p_memory_requirements MemoryRequirements)

pub type PFN_vkGetBufferMemoryRequirements = fn (device Device, buffer Buffer, mut p_memory_requirements MemoryRequirements)

@[inline]
pub fn get_buffer_memory_requirements(device Device,
	buffer Buffer,
	mut p_memory_requirements MemoryRequirements) {
	C.vkGetBufferMemoryRequirements(device, buffer, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetImageMemoryRequirements(device Device, image Image, mut p_memory_requirements MemoryRequirements)

pub type PFN_vkGetImageMemoryRequirements = fn (device Device, image Image, mut p_memory_requirements MemoryRequirements)

@[inline]
pub fn get_image_memory_requirements(device Device,
	image Image,
	mut p_memory_requirements MemoryRequirements) {
	C.vkGetImageMemoryRequirements(device, image, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetImageSparseMemoryRequirements(device Device, image Image, p_sparse_memory_requirement_count &u32, mut p_sparse_memory_requirements SparseImageMemoryRequirements)

pub type PFN_vkGetImageSparseMemoryRequirements = fn (device Device, image Image, p_sparse_memory_requirement_count &u32, mut p_sparse_memory_requirements SparseImageMemoryRequirements)

@[inline]
pub fn get_image_sparse_memory_requirements(device Device,
	image Image,
	p_sparse_memory_requirement_count &u32,
	mut p_sparse_memory_requirements SparseImageMemoryRequirements) {
	C.vkGetImageSparseMemoryRequirements(device, image, p_sparse_memory_requirement_count, mut
		p_sparse_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceSparseImageFormatProperties(physical_device PhysicalDevice, format Format, type_param ImageType, samples SampleCountFlagBits, usage ImageUsageFlags, tiling ImageTiling, p_property_count &u32, mut p_properties SparseImageFormatProperties)

pub type PFN_vkGetPhysicalDeviceSparseImageFormatProperties = fn (physical_device PhysicalDevice, format Format, type_param ImageType, samples SampleCountFlagBits, usage ImageUsageFlags, tiling ImageTiling, p_property_count &u32, mut p_properties SparseImageFormatProperties)

@[inline]
pub fn get_physical_device_sparse_image_format_properties(physical_device PhysicalDevice,
	format Format,
	type_param ImageType,
	samples SampleCountFlagBits,
	usage ImageUsageFlags,
	tiling ImageTiling,
	p_property_count &u32,
	mut p_properties SparseImageFormatProperties) {
	C.vkGetPhysicalDeviceSparseImageFormatProperties(physical_device, format, type_param,
		samples, usage, tiling, p_property_count, mut p_properties)
}

@[keep_args_alive]
fn C.vkQueueBindSparse(queue Queue, bind_info_count u32, p_bind_info &BindSparseInfo, fence Fence) Result

pub type PFN_vkQueueBindSparse = fn (queue Queue, bind_info_count u32, p_bind_info &BindSparseInfo, fence Fence) Result

@[inline]
pub fn queue_bind_sparse(queue Queue,
	bind_info_count u32,
	p_bind_info &BindSparseInfo,
	fence Fence) Result {
	return C.vkQueueBindSparse(queue, bind_info_count, p_bind_info, fence)
}

@[keep_args_alive]
fn C.vkCreateFence(device Device, p_create_info &FenceCreateInfo, p_allocator &AllocationCallbacks, p_fence &Fence) Result

pub type PFN_vkCreateFence = fn (device Device, p_create_info &FenceCreateInfo, p_allocator &AllocationCallbacks, p_fence &Fence) Result

@[inline]
pub fn create_fence(device Device,
	p_create_info &FenceCreateInfo,
	p_allocator &AllocationCallbacks,
	p_fence &Fence) Result {
	return C.vkCreateFence(device, p_create_info, p_allocator, p_fence)
}

@[keep_args_alive]
fn C.vkDestroyFence(device Device, fence Fence, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyFence = fn (device Device, fence Fence, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_fence(device Device,
	fence Fence,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyFence(device, fence, p_allocator)
}

@[keep_args_alive]
fn C.vkResetFences(device Device, fence_count u32, p_fences &Fence) Result

pub type PFN_vkResetFences = fn (device Device, fence_count u32, p_fences &Fence) Result

@[inline]
pub fn reset_fences(device Device,
	fence_count u32,
	p_fences &Fence) Result {
	return C.vkResetFences(device, fence_count, p_fences)
}

@[keep_args_alive]
fn C.vkGetFenceStatus(device Device, fence Fence) Result

pub type PFN_vkGetFenceStatus = fn (device Device, fence Fence) Result

@[inline]
pub fn get_fence_status(device Device,
	fence Fence) Result {
	return C.vkGetFenceStatus(device, fence)
}

@[keep_args_alive]
fn C.vkWaitForFences(device Device, fence_count u32, p_fences &Fence, wait_all Bool32, timeout u64) Result

pub type PFN_vkWaitForFences = fn (device Device, fence_count u32, p_fences &Fence, wait_all Bool32, timeout u64) Result

@[inline]
pub fn wait_for_fences(device Device,
	fence_count u32,
	p_fences &Fence,
	wait_all Bool32,
	timeout u64) Result {
	return C.vkWaitForFences(device, fence_count, p_fences, wait_all, timeout)
}

@[keep_args_alive]
fn C.vkCreateSemaphore(device Device, p_create_info &SemaphoreCreateInfo, p_allocator &AllocationCallbacks, p_semaphore &Semaphore) Result

pub type PFN_vkCreateSemaphore = fn (device Device, p_create_info &SemaphoreCreateInfo, p_allocator &AllocationCallbacks, p_semaphore &Semaphore) Result

@[inline]
pub fn create_semaphore(device Device,
	p_create_info &SemaphoreCreateInfo,
	p_allocator &AllocationCallbacks,
	p_semaphore &Semaphore) Result {
	return C.vkCreateSemaphore(device, p_create_info, p_allocator, p_semaphore)
}

@[keep_args_alive]
fn C.vkDestroySemaphore(device Device, semaphore Semaphore, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroySemaphore = fn (device Device, semaphore Semaphore, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_semaphore(device Device,
	semaphore Semaphore,
	p_allocator &AllocationCallbacks) {
	C.vkDestroySemaphore(device, semaphore, p_allocator)
}

@[keep_args_alive]
fn C.vkCreateQueryPool(device Device, p_create_info &QueryPoolCreateInfo, p_allocator &AllocationCallbacks, p_query_pool &QueryPool) Result

pub type PFN_vkCreateQueryPool = fn (device Device, p_create_info &QueryPoolCreateInfo, p_allocator &AllocationCallbacks, p_query_pool &QueryPool) Result

@[inline]
pub fn create_query_pool(device Device,
	p_create_info &QueryPoolCreateInfo,
	p_allocator &AllocationCallbacks,
	p_query_pool &QueryPool) Result {
	return C.vkCreateQueryPool(device, p_create_info, p_allocator, p_query_pool)
}

@[keep_args_alive]
fn C.vkDestroyQueryPool(device Device, query_pool QueryPool, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyQueryPool = fn (device Device, query_pool QueryPool, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_query_pool(device Device,
	query_pool QueryPool,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyQueryPool(device, query_pool, p_allocator)
}

@[keep_args_alive]
fn C.vkGetQueryPoolResults(device Device, query_pool QueryPool, first_query u32, query_count u32, data_size usize, p_data voidptr, stride DeviceSize, flags QueryResultFlags) Result

pub type PFN_vkGetQueryPoolResults = fn (device Device, query_pool QueryPool, first_query u32, query_count u32, data_size usize, p_data voidptr, stride DeviceSize, flags QueryResultFlags) Result

@[inline]
pub fn get_query_pool_results(device Device,
	query_pool QueryPool,
	first_query u32,
	query_count u32,
	data_size usize,
	p_data voidptr,
	stride DeviceSize,
	flags QueryResultFlags) Result {
	return C.vkGetQueryPoolResults(device, query_pool, first_query, query_count, data_size,
		p_data, stride, flags)
}

@[keep_args_alive]
fn C.vkCreateBuffer(device Device, p_create_info &BufferCreateInfo, p_allocator &AllocationCallbacks, p_buffer &Buffer) Result

pub type PFN_vkCreateBuffer = fn (device Device, p_create_info &BufferCreateInfo, p_allocator &AllocationCallbacks, p_buffer &Buffer) Result

@[inline]
pub fn create_buffer(device Device,
	p_create_info &BufferCreateInfo,
	p_allocator &AllocationCallbacks,
	p_buffer &Buffer) Result {
	return C.vkCreateBuffer(device, p_create_info, p_allocator, p_buffer)
}

@[keep_args_alive]
fn C.vkDestroyBuffer(device Device, buffer Buffer, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyBuffer = fn (device Device, buffer Buffer, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_buffer(device Device,
	buffer Buffer,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyBuffer(device, buffer, p_allocator)
}

@[keep_args_alive]
fn C.vkCreateImage(device Device, p_create_info &ImageCreateInfo, p_allocator &AllocationCallbacks, p_image &Image) Result

pub type PFN_vkCreateImage = fn (device Device, p_create_info &ImageCreateInfo, p_allocator &AllocationCallbacks, p_image &Image) Result

@[inline]
pub fn create_image(device Device,
	p_create_info &ImageCreateInfo,
	p_allocator &AllocationCallbacks,
	p_image &Image) Result {
	return C.vkCreateImage(device, p_create_info, p_allocator, p_image)
}

@[keep_args_alive]
fn C.vkDestroyImage(device Device, image Image, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyImage = fn (device Device, image Image, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_image(device Device,
	image Image,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyImage(device, image, p_allocator)
}

@[keep_args_alive]
fn C.vkGetImageSubresourceLayout(device Device, image Image, p_subresource &ImageSubresource, mut p_layout SubresourceLayout)

pub type PFN_vkGetImageSubresourceLayout = fn (device Device, image Image, p_subresource &ImageSubresource, mut p_layout SubresourceLayout)

@[inline]
pub fn get_image_subresource_layout(device Device,
	image Image,
	p_subresource &ImageSubresource,
	mut p_layout SubresourceLayout) {
	C.vkGetImageSubresourceLayout(device, image, p_subresource, mut p_layout)
}

@[keep_args_alive]
fn C.vkCreateImageView(device Device, p_create_info &ImageViewCreateInfo, p_allocator &AllocationCallbacks, p_view &ImageView) Result

pub type PFN_vkCreateImageView = fn (device Device, p_create_info &ImageViewCreateInfo, p_allocator &AllocationCallbacks, p_view &ImageView) Result

@[inline]
pub fn create_image_view(device Device,
	p_create_info &ImageViewCreateInfo,
	p_allocator &AllocationCallbacks,
	p_view &ImageView) Result {
	return C.vkCreateImageView(device, p_create_info, p_allocator, p_view)
}

@[keep_args_alive]
fn C.vkDestroyImageView(device Device, image_view ImageView, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyImageView = fn (device Device, image_view ImageView, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_image_view(device Device,
	image_view ImageView,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyImageView(device, image_view, p_allocator)
}

@[keep_args_alive]
fn C.vkCreateCommandPool(device Device, p_create_info &CommandPoolCreateInfo, p_allocator &AllocationCallbacks, p_command_pool &CommandPool) Result

pub type PFN_vkCreateCommandPool = fn (device Device, p_create_info &CommandPoolCreateInfo, p_allocator &AllocationCallbacks, p_command_pool &CommandPool) Result

@[inline]
pub fn create_command_pool(device Device,
	p_create_info &CommandPoolCreateInfo,
	p_allocator &AllocationCallbacks,
	p_command_pool &CommandPool) Result {
	return C.vkCreateCommandPool(device, p_create_info, p_allocator, p_command_pool)
}

@[keep_args_alive]
fn C.vkDestroyCommandPool(device Device, command_pool CommandPool, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyCommandPool = fn (device Device, command_pool CommandPool, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_command_pool(device Device,
	command_pool CommandPool,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyCommandPool(device, command_pool, p_allocator)
}

@[keep_args_alive]
fn C.vkResetCommandPool(device Device, command_pool CommandPool, flags CommandPoolResetFlags) Result

pub type PFN_vkResetCommandPool = fn (device Device, command_pool CommandPool, flags CommandPoolResetFlags) Result

@[inline]
pub fn reset_command_pool(device Device,
	command_pool CommandPool,
	flags CommandPoolResetFlags) Result {
	return C.vkResetCommandPool(device, command_pool, flags)
}

@[keep_args_alive]
fn C.vkAllocateCommandBuffers(device Device, p_allocate_info &CommandBufferAllocateInfo, p_command_buffers &CommandBuffer) Result

pub type PFN_vkAllocateCommandBuffers = fn (device Device, p_allocate_info &CommandBufferAllocateInfo, p_command_buffers &CommandBuffer) Result

@[inline]
pub fn allocate_command_buffers(device Device,
	p_allocate_info &CommandBufferAllocateInfo,
	p_command_buffers &CommandBuffer) Result {
	return C.vkAllocateCommandBuffers(device, p_allocate_info, p_command_buffers)
}

@[keep_args_alive]
fn C.vkFreeCommandBuffers(device Device, command_pool CommandPool, command_buffer_count u32, p_command_buffers &CommandBuffer)

pub type PFN_vkFreeCommandBuffers = fn (device Device, command_pool CommandPool, command_buffer_count u32, p_command_buffers &CommandBuffer)

@[inline]
pub fn free_command_buffers(device Device,
	command_pool CommandPool,
	command_buffer_count u32,
	p_command_buffers &CommandBuffer) {
	C.vkFreeCommandBuffers(device, command_pool, command_buffer_count, p_command_buffers)
}

@[keep_args_alive]
fn C.vkBeginCommandBuffer(command_buffer CommandBuffer, p_begin_info &CommandBufferBeginInfo) Result

pub type PFN_vkBeginCommandBuffer = fn (command_buffer CommandBuffer, p_begin_info &CommandBufferBeginInfo) Result

@[inline]
pub fn begin_command_buffer(command_buffer CommandBuffer,
	p_begin_info &CommandBufferBeginInfo) Result {
	return C.vkBeginCommandBuffer(command_buffer, p_begin_info)
}

@[keep_args_alive]
fn C.vkEndCommandBuffer(command_buffer CommandBuffer) Result

pub type PFN_vkEndCommandBuffer = fn (command_buffer CommandBuffer) Result

@[inline]
pub fn end_command_buffer(command_buffer CommandBuffer) Result {
	return C.vkEndCommandBuffer(command_buffer)
}

@[keep_args_alive]
fn C.vkResetCommandBuffer(command_buffer CommandBuffer, flags CommandBufferResetFlags) Result

pub type PFN_vkResetCommandBuffer = fn (command_buffer CommandBuffer, flags CommandBufferResetFlags) Result

@[inline]
pub fn reset_command_buffer(command_buffer CommandBuffer,
	flags CommandBufferResetFlags) Result {
	return C.vkResetCommandBuffer(command_buffer, flags)
}

@[keep_args_alive]
fn C.vkCmdCopyBuffer(command_buffer CommandBuffer, src_buffer Buffer, dst_buffer Buffer, region_count u32, p_regions &BufferCopy)

pub type PFN_vkCmdCopyBuffer = fn (command_buffer CommandBuffer, src_buffer Buffer, dst_buffer Buffer, region_count u32, p_regions &BufferCopy)

@[inline]
pub fn cmd_copy_buffer(command_buffer CommandBuffer,
	src_buffer Buffer,
	dst_buffer Buffer,
	region_count u32,
	p_regions &BufferCopy) {
	C.vkCmdCopyBuffer(command_buffer, src_buffer, dst_buffer, region_count, p_regions)
}

@[keep_args_alive]
fn C.vkCmdCopyImage(command_buffer CommandBuffer, src_image Image, src_image_layout ImageLayout, dst_image Image, dst_image_layout ImageLayout, region_count u32, p_regions &ImageCopy)

pub type PFN_vkCmdCopyImage = fn (command_buffer CommandBuffer, src_image Image, src_image_layout ImageLayout, dst_image Image, dst_image_layout ImageLayout, region_count u32, p_regions &ImageCopy)

@[inline]
pub fn cmd_copy_image(command_buffer CommandBuffer,
	src_image Image,
	src_image_layout ImageLayout,
	dst_image Image,
	dst_image_layout ImageLayout,
	region_count u32,
	p_regions &ImageCopy) {
	C.vkCmdCopyImage(command_buffer, src_image, src_image_layout, dst_image, dst_image_layout,
		region_count, p_regions)
}

@[keep_args_alive]
fn C.vkCmdCopyBufferToImage(command_buffer CommandBuffer, src_buffer Buffer, dst_image Image, dst_image_layout ImageLayout, region_count u32, p_regions &BufferImageCopy)

pub type PFN_vkCmdCopyBufferToImage = fn (command_buffer CommandBuffer, src_buffer Buffer, dst_image Image, dst_image_layout ImageLayout, region_count u32, p_regions &BufferImageCopy)

@[inline]
pub fn cmd_copy_buffer_to_image(command_buffer CommandBuffer,
	src_buffer Buffer,
	dst_image Image,
	dst_image_layout ImageLayout,
	region_count u32,
	p_regions &BufferImageCopy) {
	C.vkCmdCopyBufferToImage(command_buffer, src_buffer, dst_image, dst_image_layout,
		region_count, p_regions)
}

@[keep_args_alive]
fn C.vkCmdCopyImageToBuffer(command_buffer CommandBuffer, src_image Image, src_image_layout ImageLayout, dst_buffer Buffer, region_count u32, p_regions &BufferImageCopy)

pub type PFN_vkCmdCopyImageToBuffer = fn (command_buffer CommandBuffer, src_image Image, src_image_layout ImageLayout, dst_buffer Buffer, region_count u32, p_regions &BufferImageCopy)

@[inline]
pub fn cmd_copy_image_to_buffer(command_buffer CommandBuffer,
	src_image Image,
	src_image_layout ImageLayout,
	dst_buffer Buffer,
	region_count u32,
	p_regions &BufferImageCopy) {
	C.vkCmdCopyImageToBuffer(command_buffer, src_image, src_image_layout, dst_buffer,
		region_count, p_regions)
}

@[keep_args_alive]
fn C.vkCmdUpdateBuffer(command_buffer CommandBuffer, dst_buffer Buffer, dst_offset DeviceSize, data_size DeviceSize, p_data voidptr)

pub type PFN_vkCmdUpdateBuffer = fn (command_buffer CommandBuffer, dst_buffer Buffer, dst_offset DeviceSize, data_size DeviceSize, p_data voidptr)

@[inline]
pub fn cmd_update_buffer(command_buffer CommandBuffer,
	dst_buffer Buffer,
	dst_offset DeviceSize,
	data_size DeviceSize,
	p_data voidptr) {
	C.vkCmdUpdateBuffer(command_buffer, dst_buffer, dst_offset, data_size, p_data)
}

@[keep_args_alive]
fn C.vkCmdFillBuffer(command_buffer CommandBuffer, dst_buffer Buffer, dst_offset DeviceSize, size DeviceSize, data u32)

pub type PFN_vkCmdFillBuffer = fn (command_buffer CommandBuffer, dst_buffer Buffer, dst_offset DeviceSize, size DeviceSize, data u32)

@[inline]
pub fn cmd_fill_buffer(command_buffer CommandBuffer,
	dst_buffer Buffer,
	dst_offset DeviceSize,
	size DeviceSize,
	data u32) {
	C.vkCmdFillBuffer(command_buffer, dst_buffer, dst_offset, size, data)
}

@[keep_args_alive]
fn C.vkCmdPipelineBarrier(command_buffer CommandBuffer, src_stage_mask PipelineStageFlags, dst_stage_mask PipelineStageFlags, dependency_flags DependencyFlags, memory_barrier_count u32, p_memory_barriers &MemoryBarrier, buffer_memory_barrier_count u32, p_buffer_memory_barriers &BufferMemoryBarrier, image_memory_barrier_count u32, p_image_memory_barriers &ImageMemoryBarrier)

pub type PFN_vkCmdPipelineBarrier = fn (command_buffer CommandBuffer, src_stage_mask PipelineStageFlags, dst_stage_mask PipelineStageFlags, dependency_flags DependencyFlags, memory_barrier_count u32, p_memory_barriers &MemoryBarrier, buffer_memory_barrier_count u32, p_buffer_memory_barriers &BufferMemoryBarrier, image_memory_barrier_count u32, p_image_memory_barriers &ImageMemoryBarrier)

@[inline]
pub fn cmd_pipeline_barrier(command_buffer CommandBuffer,
	src_stage_mask PipelineStageFlags,
	dst_stage_mask PipelineStageFlags,
	dependency_flags DependencyFlags,
	memory_barrier_count u32,
	p_memory_barriers &MemoryBarrier,
	buffer_memory_barrier_count u32,
	p_buffer_memory_barriers &BufferMemoryBarrier,
	image_memory_barrier_count u32,
	p_image_memory_barriers &ImageMemoryBarrier) {
	C.vkCmdPipelineBarrier(command_buffer, src_stage_mask, dst_stage_mask, dependency_flags,
		memory_barrier_count, p_memory_barriers, buffer_memory_barrier_count, p_buffer_memory_barriers,
		image_memory_barrier_count, p_image_memory_barriers)
}

@[keep_args_alive]
fn C.vkCmdBeginQuery(command_buffer CommandBuffer, query_pool QueryPool, query u32, flags QueryControlFlags)

pub type PFN_vkCmdBeginQuery = fn (command_buffer CommandBuffer, query_pool QueryPool, query u32, flags QueryControlFlags)

@[inline]
pub fn cmd_begin_query(command_buffer CommandBuffer,
	query_pool QueryPool,
	query u32,
	flags QueryControlFlags) {
	C.vkCmdBeginQuery(command_buffer, query_pool, query, flags)
}

@[keep_args_alive]
fn C.vkCmdEndQuery(command_buffer CommandBuffer, query_pool QueryPool, query u32)

pub type PFN_vkCmdEndQuery = fn (command_buffer CommandBuffer, query_pool QueryPool, query u32)

@[inline]
pub fn cmd_end_query(command_buffer CommandBuffer,
	query_pool QueryPool,
	query u32) {
	C.vkCmdEndQuery(command_buffer, query_pool, query)
}

@[keep_args_alive]
fn C.vkCmdResetQueryPool(command_buffer CommandBuffer, query_pool QueryPool, first_query u32, query_count u32)

pub type PFN_vkCmdResetQueryPool = fn (command_buffer CommandBuffer, query_pool QueryPool, first_query u32, query_count u32)

@[inline]
pub fn cmd_reset_query_pool(command_buffer CommandBuffer,
	query_pool QueryPool,
	first_query u32,
	query_count u32) {
	C.vkCmdResetQueryPool(command_buffer, query_pool, first_query, query_count)
}

@[keep_args_alive]
fn C.vkCmdWriteTimestamp(command_buffer CommandBuffer, pipeline_stage PipelineStageFlagBits, query_pool QueryPool, query u32)

pub type PFN_vkCmdWriteTimestamp = fn (command_buffer CommandBuffer, pipeline_stage PipelineStageFlagBits, query_pool QueryPool, query u32)

@[inline]
pub fn cmd_write_timestamp(command_buffer CommandBuffer,
	pipeline_stage PipelineStageFlagBits,
	query_pool QueryPool,
	query u32) {
	C.vkCmdWriteTimestamp(command_buffer, pipeline_stage, query_pool, query)
}

@[keep_args_alive]
fn C.vkCmdCopyQueryPoolResults(command_buffer CommandBuffer, query_pool QueryPool, first_query u32, query_count u32, dst_buffer Buffer, dst_offset DeviceSize, stride DeviceSize, flags QueryResultFlags)

pub type PFN_vkCmdCopyQueryPoolResults = fn (command_buffer CommandBuffer, query_pool QueryPool, first_query u32, query_count u32, dst_buffer Buffer, dst_offset DeviceSize, stride DeviceSize, flags QueryResultFlags)

@[inline]
pub fn cmd_copy_query_pool_results(command_buffer CommandBuffer,
	query_pool QueryPool,
	first_query u32,
	query_count u32,
	dst_buffer Buffer,
	dst_offset DeviceSize,
	stride DeviceSize,
	flags QueryResultFlags) {
	C.vkCmdCopyQueryPoolResults(command_buffer, query_pool, first_query, query_count,
		dst_buffer, dst_offset, stride, flags)
}

@[keep_args_alive]
fn C.vkCmdExecuteCommands(command_buffer CommandBuffer, command_buffer_count u32, p_command_buffers &CommandBuffer)

pub type PFN_vkCmdExecuteCommands = fn (command_buffer CommandBuffer, command_buffer_count u32, p_command_buffers &CommandBuffer)

@[inline]
pub fn cmd_execute_commands(command_buffer CommandBuffer,
	command_buffer_count u32,
	p_command_buffers &CommandBuffer) {
	C.vkCmdExecuteCommands(command_buffer, command_buffer_count, p_command_buffers)
}

@[keep_args_alive]
fn C.vkCreateEvent(device Device, p_create_info &EventCreateInfo, p_allocator &AllocationCallbacks, p_event &Event) Result

pub type PFN_vkCreateEvent = fn (device Device, p_create_info &EventCreateInfo, p_allocator &AllocationCallbacks, p_event &Event) Result

@[inline]
pub fn create_event(device Device,
	p_create_info &EventCreateInfo,
	p_allocator &AllocationCallbacks,
	p_event &Event) Result {
	return C.vkCreateEvent(device, p_create_info, p_allocator, p_event)
}

@[keep_args_alive]
fn C.vkDestroyEvent(device Device, event Event, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyEvent = fn (device Device, event Event, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_event(device Device,
	event Event,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyEvent(device, event, p_allocator)
}

@[keep_args_alive]
fn C.vkGetEventStatus(device Device, event Event) Result

pub type PFN_vkGetEventStatus = fn (device Device, event Event) Result

@[inline]
pub fn get_event_status(device Device,
	event Event) Result {
	return C.vkGetEventStatus(device, event)
}

@[keep_args_alive]
fn C.vkSetEvent(device Device, event Event) Result

pub type PFN_vkSetEvent = fn (device Device, event Event) Result

@[inline]
pub fn set_event(device Device,
	event Event) Result {
	return C.vkSetEvent(device, event)
}

@[keep_args_alive]
fn C.vkResetEvent(device Device, event Event) Result

pub type PFN_vkResetEvent = fn (device Device, event Event) Result

@[inline]
pub fn reset_event(device Device,
	event Event) Result {
	return C.vkResetEvent(device, event)
}

@[keep_args_alive]
fn C.vkCreateBufferView(device Device, p_create_info &BufferViewCreateInfo, p_allocator &AllocationCallbacks, p_view &BufferView) Result

pub type PFN_vkCreateBufferView = fn (device Device, p_create_info &BufferViewCreateInfo, p_allocator &AllocationCallbacks, p_view &BufferView) Result

@[inline]
pub fn create_buffer_view(device Device,
	p_create_info &BufferViewCreateInfo,
	p_allocator &AllocationCallbacks,
	p_view &BufferView) Result {
	return C.vkCreateBufferView(device, p_create_info, p_allocator, p_view)
}

@[keep_args_alive]
fn C.vkDestroyBufferView(device Device, buffer_view BufferView, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyBufferView = fn (device Device, buffer_view BufferView, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_buffer_view(device Device,
	buffer_view BufferView,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyBufferView(device, buffer_view, p_allocator)
}

@[keep_args_alive]
fn C.vkCreateShaderModule(device Device, p_create_info &ShaderModuleCreateInfo, p_allocator &AllocationCallbacks, p_shader_module &ShaderModule) Result

pub type PFN_vkCreateShaderModule = fn (device Device, p_create_info &ShaderModuleCreateInfo, p_allocator &AllocationCallbacks, p_shader_module &ShaderModule) Result

@[inline]
pub fn create_shader_module(device Device,
	p_create_info &ShaderModuleCreateInfo,
	p_allocator &AllocationCallbacks,
	p_shader_module &ShaderModule) Result {
	return C.vkCreateShaderModule(device, p_create_info, p_allocator, p_shader_module)
}

@[keep_args_alive]
fn C.vkDestroyShaderModule(device Device, shader_module ShaderModule, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyShaderModule = fn (device Device, shader_module ShaderModule, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_shader_module(device Device,
	shader_module ShaderModule,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyShaderModule(device, shader_module, p_allocator)
}

@[keep_args_alive]
fn C.vkCreatePipelineCache(device Device, p_create_info &PipelineCacheCreateInfo, p_allocator &AllocationCallbacks, p_pipeline_cache &PipelineCache) Result

pub type PFN_vkCreatePipelineCache = fn (device Device, p_create_info &PipelineCacheCreateInfo, p_allocator &AllocationCallbacks, p_pipeline_cache &PipelineCache) Result

@[inline]
pub fn create_pipeline_cache(device Device,
	p_create_info &PipelineCacheCreateInfo,
	p_allocator &AllocationCallbacks,
	p_pipeline_cache &PipelineCache) Result {
	return C.vkCreatePipelineCache(device, p_create_info, p_allocator, p_pipeline_cache)
}

@[keep_args_alive]
fn C.vkDestroyPipelineCache(device Device, pipeline_cache PipelineCache, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyPipelineCache = fn (device Device, pipeline_cache PipelineCache, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_pipeline_cache(device Device,
	pipeline_cache PipelineCache,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyPipelineCache(device, pipeline_cache, p_allocator)
}

@[keep_args_alive]
fn C.vkGetPipelineCacheData(device Device, pipeline_cache PipelineCache, p_data_size &usize, p_data voidptr) Result

pub type PFN_vkGetPipelineCacheData = fn (device Device, pipeline_cache PipelineCache, p_data_size &usize, p_data voidptr) Result

@[inline]
pub fn get_pipeline_cache_data(device Device,
	pipeline_cache PipelineCache,
	p_data_size &usize,
	p_data voidptr) Result {
	return C.vkGetPipelineCacheData(device, pipeline_cache, p_data_size, p_data)
}

@[keep_args_alive]
fn C.vkMergePipelineCaches(device Device, dst_cache PipelineCache, src_cache_count u32, p_src_caches &PipelineCache) Result

pub type PFN_vkMergePipelineCaches = fn (device Device, dst_cache PipelineCache, src_cache_count u32, p_src_caches &PipelineCache) Result

@[inline]
pub fn merge_pipeline_caches(device Device,
	dst_cache PipelineCache,
	src_cache_count u32,
	p_src_caches &PipelineCache) Result {
	return C.vkMergePipelineCaches(device, dst_cache, src_cache_count, p_src_caches)
}

@[keep_args_alive]
fn C.vkCreateComputePipelines(device Device, pipeline_cache PipelineCache, create_info_count u32, p_create_infos &ComputePipelineCreateInfo, p_allocator &AllocationCallbacks, p_pipelines &Pipeline) Result

pub type PFN_vkCreateComputePipelines = fn (device Device, pipeline_cache PipelineCache, create_info_count u32, p_create_infos &ComputePipelineCreateInfo, p_allocator &AllocationCallbacks, p_pipelines &Pipeline) Result

@[inline]
pub fn create_compute_pipelines(device Device,
	pipeline_cache PipelineCache,
	create_info_count u32,
	p_create_infos &ComputePipelineCreateInfo,
	p_allocator &AllocationCallbacks,
	p_pipelines &Pipeline) Result {
	return C.vkCreateComputePipelines(device, pipeline_cache, create_info_count, p_create_infos,
		p_allocator, p_pipelines)
}

@[keep_args_alive]
fn C.vkDestroyPipeline(device Device, pipeline Pipeline, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyPipeline = fn (device Device, pipeline Pipeline, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_pipeline(device Device,
	pipeline Pipeline,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyPipeline(device, pipeline, p_allocator)
}

@[keep_args_alive]
fn C.vkCreatePipelineLayout(device Device, p_create_info &PipelineLayoutCreateInfo, p_allocator &AllocationCallbacks, p_pipeline_layout &PipelineLayout) Result

pub type PFN_vkCreatePipelineLayout = fn (device Device, p_create_info &PipelineLayoutCreateInfo, p_allocator &AllocationCallbacks, p_pipeline_layout &PipelineLayout) Result

@[inline]
pub fn create_pipeline_layout(device Device,
	p_create_info &PipelineLayoutCreateInfo,
	p_allocator &AllocationCallbacks,
	p_pipeline_layout &PipelineLayout) Result {
	return C.vkCreatePipelineLayout(device, p_create_info, p_allocator, p_pipeline_layout)
}

@[keep_args_alive]
fn C.vkDestroyPipelineLayout(device Device, pipeline_layout PipelineLayout, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyPipelineLayout = fn (device Device, pipeline_layout PipelineLayout, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_pipeline_layout(device Device,
	pipeline_layout PipelineLayout,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyPipelineLayout(device, pipeline_layout, p_allocator)
}

@[keep_args_alive]
fn C.vkCreateSampler(device Device, p_create_info &SamplerCreateInfo, p_allocator &AllocationCallbacks, p_sampler &Sampler) Result

pub type PFN_vkCreateSampler = fn (device Device, p_create_info &SamplerCreateInfo, p_allocator &AllocationCallbacks, p_sampler &Sampler) Result

@[inline]
pub fn create_sampler(device Device,
	p_create_info &SamplerCreateInfo,
	p_allocator &AllocationCallbacks,
	p_sampler &Sampler) Result {
	return C.vkCreateSampler(device, p_create_info, p_allocator, p_sampler)
}

@[keep_args_alive]
fn C.vkDestroySampler(device Device, sampler Sampler, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroySampler = fn (device Device, sampler Sampler, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_sampler(device Device,
	sampler Sampler,
	p_allocator &AllocationCallbacks) {
	C.vkDestroySampler(device, sampler, p_allocator)
}

@[keep_args_alive]
fn C.vkCreateDescriptorSetLayout(device Device, p_create_info &DescriptorSetLayoutCreateInfo, p_allocator &AllocationCallbacks, p_set_layout &DescriptorSetLayout) Result

pub type PFN_vkCreateDescriptorSetLayout = fn (device Device, p_create_info &DescriptorSetLayoutCreateInfo, p_allocator &AllocationCallbacks, p_set_layout &DescriptorSetLayout) Result

@[inline]
pub fn create_descriptor_set_layout(device Device,
	p_create_info &DescriptorSetLayoutCreateInfo,
	p_allocator &AllocationCallbacks,
	p_set_layout &DescriptorSetLayout) Result {
	return C.vkCreateDescriptorSetLayout(device, p_create_info, p_allocator, p_set_layout)
}

@[keep_args_alive]
fn C.vkDestroyDescriptorSetLayout(device Device, descriptor_set_layout DescriptorSetLayout, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyDescriptorSetLayout = fn (device Device, descriptor_set_layout DescriptorSetLayout, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_descriptor_set_layout(device Device,
	descriptor_set_layout DescriptorSetLayout,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyDescriptorSetLayout(device, descriptor_set_layout, p_allocator)
}

@[keep_args_alive]
fn C.vkCreateDescriptorPool(device Device, p_create_info &DescriptorPoolCreateInfo, p_allocator &AllocationCallbacks, p_descriptor_pool &DescriptorPool) Result

pub type PFN_vkCreateDescriptorPool = fn (device Device, p_create_info &DescriptorPoolCreateInfo, p_allocator &AllocationCallbacks, p_descriptor_pool &DescriptorPool) Result

@[inline]
pub fn create_descriptor_pool(device Device,
	p_create_info &DescriptorPoolCreateInfo,
	p_allocator &AllocationCallbacks,
	p_descriptor_pool &DescriptorPool) Result {
	return C.vkCreateDescriptorPool(device, p_create_info, p_allocator, p_descriptor_pool)
}

@[keep_args_alive]
fn C.vkDestroyDescriptorPool(device Device, descriptor_pool DescriptorPool, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyDescriptorPool = fn (device Device, descriptor_pool DescriptorPool, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_descriptor_pool(device Device,
	descriptor_pool DescriptorPool,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyDescriptorPool(device, descriptor_pool, p_allocator)
}

@[keep_args_alive]
fn C.vkResetDescriptorPool(device Device, descriptor_pool DescriptorPool, flags DescriptorPoolResetFlags) Result

pub type PFN_vkResetDescriptorPool = fn (device Device, descriptor_pool DescriptorPool, flags DescriptorPoolResetFlags) Result

@[inline]
pub fn reset_descriptor_pool(device Device,
	descriptor_pool DescriptorPool,
	flags DescriptorPoolResetFlags) Result {
	return C.vkResetDescriptorPool(device, descriptor_pool, flags)
}

@[keep_args_alive]
fn C.vkAllocateDescriptorSets(device Device, p_allocate_info &DescriptorSetAllocateInfo, p_descriptor_sets &DescriptorSet) Result

pub type PFN_vkAllocateDescriptorSets = fn (device Device, p_allocate_info &DescriptorSetAllocateInfo, p_descriptor_sets &DescriptorSet) Result

@[inline]
pub fn allocate_descriptor_sets(device Device,
	p_allocate_info &DescriptorSetAllocateInfo,
	p_descriptor_sets &DescriptorSet) Result {
	return C.vkAllocateDescriptorSets(device, p_allocate_info, p_descriptor_sets)
}

@[keep_args_alive]
fn C.vkFreeDescriptorSets(device Device, descriptor_pool DescriptorPool, descriptor_set_count u32, p_descriptor_sets &DescriptorSet) Result

pub type PFN_vkFreeDescriptorSets = fn (device Device, descriptor_pool DescriptorPool, descriptor_set_count u32, p_descriptor_sets &DescriptorSet) Result

@[inline]
pub fn free_descriptor_sets(device Device,
	descriptor_pool DescriptorPool,
	descriptor_set_count u32,
	p_descriptor_sets &DescriptorSet) Result {
	return C.vkFreeDescriptorSets(device, descriptor_pool, descriptor_set_count, p_descriptor_sets)
}

@[keep_args_alive]
fn C.vkUpdateDescriptorSets(device Device, descriptor_write_count u32, p_descriptor_writes &WriteDescriptorSet, descriptor_copy_count u32, p_descriptor_copies &CopyDescriptorSet)

pub type PFN_vkUpdateDescriptorSets = fn (device Device, descriptor_write_count u32, p_descriptor_writes &WriteDescriptorSet, descriptor_copy_count u32, p_descriptor_copies &CopyDescriptorSet)

@[inline]
pub fn update_descriptor_sets(device Device,
	descriptor_write_count u32,
	p_descriptor_writes &WriteDescriptorSet,
	descriptor_copy_count u32,
	p_descriptor_copies &CopyDescriptorSet) {
	C.vkUpdateDescriptorSets(device, descriptor_write_count, p_descriptor_writes, descriptor_copy_count,
		p_descriptor_copies)
}

@[keep_args_alive]
fn C.vkCmdBindPipeline(command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, pipeline Pipeline)

pub type PFN_vkCmdBindPipeline = fn (command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, pipeline Pipeline)

@[inline]
pub fn cmd_bind_pipeline(command_buffer CommandBuffer,
	pipeline_bind_point PipelineBindPoint,
	pipeline Pipeline) {
	C.vkCmdBindPipeline(command_buffer, pipeline_bind_point, pipeline)
}

@[keep_args_alive]
fn C.vkCmdBindDescriptorSets(command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, layout PipelineLayout, first_set u32, descriptor_set_count u32, p_descriptor_sets &DescriptorSet, dynamic_offset_count u32, p_dynamic_offsets &u32)

pub type PFN_vkCmdBindDescriptorSets = fn (command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, layout PipelineLayout, first_set u32, descriptor_set_count u32, p_descriptor_sets &DescriptorSet, dynamic_offset_count u32, p_dynamic_offsets &u32)

@[inline]
pub fn cmd_bind_descriptor_sets(command_buffer CommandBuffer,
	pipeline_bind_point PipelineBindPoint,
	layout PipelineLayout,
	first_set u32,
	descriptor_set_count u32,
	p_descriptor_sets &DescriptorSet,
	dynamic_offset_count u32,
	p_dynamic_offsets &u32) {
	C.vkCmdBindDescriptorSets(command_buffer, pipeline_bind_point, layout, first_set,
		descriptor_set_count, p_descriptor_sets, dynamic_offset_count, p_dynamic_offsets)
}

@[keep_args_alive]
fn C.vkCmdClearColorImage(command_buffer CommandBuffer, image Image, image_layout ImageLayout, p_color &ClearColorValue, range_count u32, p_ranges &ImageSubresourceRange)

pub type PFN_vkCmdClearColorImage = fn (command_buffer CommandBuffer, image Image, image_layout ImageLayout, p_color &ClearColorValue, range_count u32, p_ranges &ImageSubresourceRange)

@[inline]
pub fn cmd_clear_color_image(command_buffer CommandBuffer,
	image Image,
	image_layout ImageLayout,
	p_color &ClearColorValue,
	range_count u32,
	p_ranges &ImageSubresourceRange) {
	C.vkCmdClearColorImage(command_buffer, image, image_layout, p_color, range_count,
		p_ranges)
}

@[keep_args_alive]
fn C.vkCmdDispatch(command_buffer CommandBuffer, group_count_x u32, group_count_y u32, group_count_z u32)

pub type PFN_vkCmdDispatch = fn (command_buffer CommandBuffer, group_count_x u32, group_count_y u32, group_count_z u32)

@[inline]
pub fn cmd_dispatch(command_buffer CommandBuffer,
	group_count_x u32,
	group_count_y u32,
	group_count_z u32) {
	C.vkCmdDispatch(command_buffer, group_count_x, group_count_y, group_count_z)
}

@[keep_args_alive]
fn C.vkCmdDispatchIndirect(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize)

pub type PFN_vkCmdDispatchIndirect = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize)

@[inline]
pub fn cmd_dispatch_indirect(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize) {
	C.vkCmdDispatchIndirect(command_buffer, buffer, offset)
}

@[keep_args_alive]
fn C.vkCmdSetEvent(command_buffer CommandBuffer, event Event, stage_mask PipelineStageFlags)

pub type PFN_vkCmdSetEvent = fn (command_buffer CommandBuffer, event Event, stage_mask PipelineStageFlags)

@[inline]
pub fn cmd_set_event(command_buffer CommandBuffer,
	event Event,
	stage_mask PipelineStageFlags) {
	C.vkCmdSetEvent(command_buffer, event, stage_mask)
}

@[keep_args_alive]
fn C.vkCmdResetEvent(command_buffer CommandBuffer, event Event, stage_mask PipelineStageFlags)

pub type PFN_vkCmdResetEvent = fn (command_buffer CommandBuffer, event Event, stage_mask PipelineStageFlags)

@[inline]
pub fn cmd_reset_event(command_buffer CommandBuffer,
	event Event,
	stage_mask PipelineStageFlags) {
	C.vkCmdResetEvent(command_buffer, event, stage_mask)
}

@[keep_args_alive]
fn C.vkCmdWaitEvents(command_buffer CommandBuffer, event_count u32, p_events &Event, src_stage_mask PipelineStageFlags, dst_stage_mask PipelineStageFlags, memory_barrier_count u32, p_memory_barriers &MemoryBarrier, buffer_memory_barrier_count u32, p_buffer_memory_barriers &BufferMemoryBarrier, image_memory_barrier_count u32, p_image_memory_barriers &ImageMemoryBarrier)

pub type PFN_vkCmdWaitEvents = fn (command_buffer CommandBuffer, event_count u32, p_events &Event, src_stage_mask PipelineStageFlags, dst_stage_mask PipelineStageFlags, memory_barrier_count u32, p_memory_barriers &MemoryBarrier, buffer_memory_barrier_count u32, p_buffer_memory_barriers &BufferMemoryBarrier, image_memory_barrier_count u32, p_image_memory_barriers &ImageMemoryBarrier)

@[inline]
pub fn cmd_wait_events(command_buffer CommandBuffer,
	event_count u32,
	p_events &Event,
	src_stage_mask PipelineStageFlags,
	dst_stage_mask PipelineStageFlags,
	memory_barrier_count u32,
	p_memory_barriers &MemoryBarrier,
	buffer_memory_barrier_count u32,
	p_buffer_memory_barriers &BufferMemoryBarrier,
	image_memory_barrier_count u32,
	p_image_memory_barriers &ImageMemoryBarrier) {
	C.vkCmdWaitEvents(command_buffer, event_count, p_events, src_stage_mask, dst_stage_mask,
		memory_barrier_count, p_memory_barriers, buffer_memory_barrier_count, p_buffer_memory_barriers,
		image_memory_barrier_count, p_image_memory_barriers)
}

@[keep_args_alive]
fn C.vkCmdPushConstants(command_buffer CommandBuffer, layout PipelineLayout, stage_flags ShaderStageFlags, offset u32, size u32, p_values voidptr)

pub type PFN_vkCmdPushConstants = fn (command_buffer CommandBuffer, layout PipelineLayout, stage_flags ShaderStageFlags, offset u32, size u32, p_values voidptr)

@[inline]
pub fn cmd_push_constants(command_buffer CommandBuffer,
	layout PipelineLayout,
	stage_flags ShaderStageFlags,
	offset u32,
	size u32,
	p_values voidptr) {
	C.vkCmdPushConstants(command_buffer, layout, stage_flags, offset, size, p_values)
}

@[keep_args_alive]
fn C.vkCreateGraphicsPipelines(device Device, pipeline_cache PipelineCache, create_info_count u32, p_create_infos &GraphicsPipelineCreateInfo, p_allocator &AllocationCallbacks, p_pipelines &Pipeline) Result

pub type PFN_vkCreateGraphicsPipelines = fn (device Device, pipeline_cache PipelineCache, create_info_count u32, p_create_infos &GraphicsPipelineCreateInfo, p_allocator &AllocationCallbacks, p_pipelines &Pipeline) Result

@[inline]
pub fn create_graphics_pipelines(device Device,
	pipeline_cache PipelineCache,
	create_info_count u32,
	p_create_infos &GraphicsPipelineCreateInfo,
	p_allocator &AllocationCallbacks,
	p_pipelines &Pipeline) Result {
	return C.vkCreateGraphicsPipelines(device, pipeline_cache, create_info_count, p_create_infos,
		p_allocator, p_pipelines)
}

@[keep_args_alive]
fn C.vkCreateFramebuffer(device Device, p_create_info &FramebufferCreateInfo, p_allocator &AllocationCallbacks, p_framebuffer &Framebuffer) Result

pub type PFN_vkCreateFramebuffer = fn (device Device, p_create_info &FramebufferCreateInfo, p_allocator &AllocationCallbacks, p_framebuffer &Framebuffer) Result

@[inline]
pub fn create_framebuffer(device Device,
	p_create_info &FramebufferCreateInfo,
	p_allocator &AllocationCallbacks,
	p_framebuffer &Framebuffer) Result {
	return C.vkCreateFramebuffer(device, p_create_info, p_allocator, p_framebuffer)
}

@[keep_args_alive]
fn C.vkDestroyFramebuffer(device Device, framebuffer Framebuffer, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyFramebuffer = fn (device Device, framebuffer Framebuffer, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_framebuffer(device Device,
	framebuffer Framebuffer,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyFramebuffer(device, framebuffer, p_allocator)
}

@[keep_args_alive]
fn C.vkCreateRenderPass(device Device, p_create_info &RenderPassCreateInfo, p_allocator &AllocationCallbacks, p_render_pass &RenderPass) Result

pub type PFN_vkCreateRenderPass = fn (device Device, p_create_info &RenderPassCreateInfo, p_allocator &AllocationCallbacks, p_render_pass &RenderPass) Result

@[inline]
pub fn create_render_pass(device Device,
	p_create_info &RenderPassCreateInfo,
	p_allocator &AllocationCallbacks,
	p_render_pass &RenderPass) Result {
	return C.vkCreateRenderPass(device, p_create_info, p_allocator, p_render_pass)
}

@[keep_args_alive]
fn C.vkDestroyRenderPass(device Device, render_pass RenderPass, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyRenderPass = fn (device Device, render_pass RenderPass, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_render_pass(device Device,
	render_pass RenderPass,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyRenderPass(device, render_pass, p_allocator)
}

@[keep_args_alive]
fn C.vkGetRenderAreaGranularity(device Device, render_pass RenderPass, mut p_granularity Extent2D)

pub type PFN_vkGetRenderAreaGranularity = fn (device Device, render_pass RenderPass, mut p_granularity Extent2D)

@[inline]
pub fn get_render_area_granularity(device Device,
	render_pass RenderPass,
	mut p_granularity Extent2D) {
	C.vkGetRenderAreaGranularity(device, render_pass, mut p_granularity)
}

@[keep_args_alive]
fn C.vkCmdSetViewport(command_buffer CommandBuffer, first_viewport u32, viewport_count u32, p_viewports &Viewport)

pub type PFN_vkCmdSetViewport = fn (command_buffer CommandBuffer, first_viewport u32, viewport_count u32, p_viewports &Viewport)

@[inline]
pub fn cmd_set_viewport(command_buffer CommandBuffer,
	first_viewport u32,
	viewport_count u32,
	p_viewports &Viewport) {
	C.vkCmdSetViewport(command_buffer, first_viewport, viewport_count, p_viewports)
}

@[keep_args_alive]
fn C.vkCmdSetScissor(command_buffer CommandBuffer, first_scissor u32, scissor_count u32, p_scissors &Rect2D)

pub type PFN_vkCmdSetScissor = fn (command_buffer CommandBuffer, first_scissor u32, scissor_count u32, p_scissors &Rect2D)

@[inline]
pub fn cmd_set_scissor(command_buffer CommandBuffer,
	first_scissor u32,
	scissor_count u32,
	p_scissors &Rect2D) {
	C.vkCmdSetScissor(command_buffer, first_scissor, scissor_count, p_scissors)
}

@[keep_args_alive]
fn C.vkCmdSetLineWidth(command_buffer CommandBuffer, line_width f32)

pub type PFN_vkCmdSetLineWidth = fn (command_buffer CommandBuffer, line_width f32)

@[inline]
pub fn cmd_set_line_width(command_buffer CommandBuffer,
	line_width f32) {
	C.vkCmdSetLineWidth(command_buffer, line_width)
}

@[keep_args_alive]
fn C.vkCmdSetDepthBias(command_buffer CommandBuffer, depth_bias_constant_factor f32, depth_bias_clamp f32, depth_bias_slope_factor f32)

pub type PFN_vkCmdSetDepthBias = fn (command_buffer CommandBuffer, depth_bias_constant_factor f32, depth_bias_clamp f32, depth_bias_slope_factor f32)

@[inline]
pub fn cmd_set_depth_bias(command_buffer CommandBuffer,
	depth_bias_constant_factor f32,
	depth_bias_clamp f32,
	depth_bias_slope_factor f32) {
	C.vkCmdSetDepthBias(command_buffer, depth_bias_constant_factor, depth_bias_clamp,
		depth_bias_slope_factor)
}

@[keep_args_alive]
fn C.vkCmdSetBlendConstants(command_buffer CommandBuffer, blend_constants [4]f32)

pub type PFN_vkCmdSetBlendConstants = fn (command_buffer CommandBuffer, blend_constants [4]f32)

@[inline]
pub fn cmd_set_blend_constants(command_buffer CommandBuffer,
	blend_constants [4]f32) {
	C.vkCmdSetBlendConstants(command_buffer, blend_constants)
}

@[keep_args_alive]
fn C.vkCmdSetDepthBounds(command_buffer CommandBuffer, min_depth_bounds f32, max_depth_bounds f32)

pub type PFN_vkCmdSetDepthBounds = fn (command_buffer CommandBuffer, min_depth_bounds f32, max_depth_bounds f32)

@[inline]
pub fn cmd_set_depth_bounds(command_buffer CommandBuffer,
	min_depth_bounds f32,
	max_depth_bounds f32) {
	C.vkCmdSetDepthBounds(command_buffer, min_depth_bounds, max_depth_bounds)
}

@[keep_args_alive]
fn C.vkCmdSetStencilCompareMask(command_buffer CommandBuffer, face_mask StencilFaceFlags, compare_mask u32)

pub type PFN_vkCmdSetStencilCompareMask = fn (command_buffer CommandBuffer, face_mask StencilFaceFlags, compare_mask u32)

@[inline]
pub fn cmd_set_stencil_compare_mask(command_buffer CommandBuffer,
	face_mask StencilFaceFlags,
	compare_mask u32) {
	C.vkCmdSetStencilCompareMask(command_buffer, face_mask, compare_mask)
}

@[keep_args_alive]
fn C.vkCmdSetStencilWriteMask(command_buffer CommandBuffer, face_mask StencilFaceFlags, write_mask u32)

pub type PFN_vkCmdSetStencilWriteMask = fn (command_buffer CommandBuffer, face_mask StencilFaceFlags, write_mask u32)

@[inline]
pub fn cmd_set_stencil_write_mask(command_buffer CommandBuffer,
	face_mask StencilFaceFlags,
	write_mask u32) {
	C.vkCmdSetStencilWriteMask(command_buffer, face_mask, write_mask)
}

@[keep_args_alive]
fn C.vkCmdSetStencilReference(command_buffer CommandBuffer, face_mask StencilFaceFlags, reference u32)

pub type PFN_vkCmdSetStencilReference = fn (command_buffer CommandBuffer, face_mask StencilFaceFlags, reference u32)

@[inline]
pub fn cmd_set_stencil_reference(command_buffer CommandBuffer,
	face_mask StencilFaceFlags,
	reference u32) {
	C.vkCmdSetStencilReference(command_buffer, face_mask, reference)
}

@[keep_args_alive]
fn C.vkCmdBindIndexBuffer(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, index_type IndexType)

pub type PFN_vkCmdBindIndexBuffer = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, index_type IndexType)

@[inline]
pub fn cmd_bind_index_buffer(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	index_type IndexType) {
	C.vkCmdBindIndexBuffer(command_buffer, buffer, offset, index_type)
}

@[keep_args_alive]
fn C.vkCmdBindVertexBuffers(command_buffer CommandBuffer, first_binding u32, binding_count u32, p_buffers &Buffer, p_offsets &DeviceSize)

pub type PFN_vkCmdBindVertexBuffers = fn (command_buffer CommandBuffer, first_binding u32, binding_count u32, p_buffers &Buffer, p_offsets &DeviceSize)

@[inline]
pub fn cmd_bind_vertex_buffers(command_buffer CommandBuffer,
	first_binding u32,
	binding_count u32,
	p_buffers &Buffer,
	p_offsets &DeviceSize) {
	C.vkCmdBindVertexBuffers(command_buffer, first_binding, binding_count, p_buffers,
		p_offsets)
}

@[keep_args_alive]
fn C.vkCmdDraw(command_buffer CommandBuffer, vertex_count u32, instance_count u32, first_vertex u32, first_instance u32)

pub type PFN_vkCmdDraw = fn (command_buffer CommandBuffer, vertex_count u32, instance_count u32, first_vertex u32, first_instance u32)

@[inline]
pub fn cmd_draw(command_buffer CommandBuffer,
	vertex_count u32,
	instance_count u32,
	first_vertex u32,
	first_instance u32) {
	C.vkCmdDraw(command_buffer, vertex_count, instance_count, first_vertex, first_instance)
}

@[keep_args_alive]
fn C.vkCmdDrawIndexed(command_buffer CommandBuffer, index_count u32, instance_count u32, first_index u32, vertex_offset i32, first_instance u32)

pub type PFN_vkCmdDrawIndexed = fn (command_buffer CommandBuffer, index_count u32, instance_count u32, first_index u32, vertex_offset i32, first_instance u32)

@[inline]
pub fn cmd_draw_indexed(command_buffer CommandBuffer,
	index_count u32,
	instance_count u32,
	first_index u32,
	vertex_offset i32,
	first_instance u32) {
	C.vkCmdDrawIndexed(command_buffer, index_count, instance_count, first_index, vertex_offset,
		first_instance)
}

@[keep_args_alive]
fn C.vkCmdDrawIndirect(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, draw_count u32, stride u32)

pub type PFN_vkCmdDrawIndirect = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_indirect(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	draw_count u32,
	stride u32) {
	C.vkCmdDrawIndirect(command_buffer, buffer, offset, draw_count, stride)
}

@[keep_args_alive]
fn C.vkCmdDrawIndexedIndirect(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, draw_count u32, stride u32)

pub type PFN_vkCmdDrawIndexedIndirect = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_indexed_indirect(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	draw_count u32,
	stride u32) {
	C.vkCmdDrawIndexedIndirect(command_buffer, buffer, offset, draw_count, stride)
}

@[keep_args_alive]
fn C.vkCmdBlitImage(command_buffer CommandBuffer, src_image Image, src_image_layout ImageLayout, dst_image Image, dst_image_layout ImageLayout, region_count u32, p_regions &ImageBlit, filter Filter)

pub type PFN_vkCmdBlitImage = fn (command_buffer CommandBuffer, src_image Image, src_image_layout ImageLayout, dst_image Image, dst_image_layout ImageLayout, region_count u32, p_regions &ImageBlit, filter Filter)

@[inline]
pub fn cmd_blit_image(command_buffer CommandBuffer,
	src_image Image,
	src_image_layout ImageLayout,
	dst_image Image,
	dst_image_layout ImageLayout,
	region_count u32,
	p_regions &ImageBlit,
	filter Filter) {
	C.vkCmdBlitImage(command_buffer, src_image, src_image_layout, dst_image, dst_image_layout,
		region_count, p_regions, filter)
}

@[keep_args_alive]
fn C.vkCmdClearDepthStencilImage(command_buffer CommandBuffer, image Image, image_layout ImageLayout, p_depth_stencil &ClearDepthStencilValue, range_count u32, p_ranges &ImageSubresourceRange)

pub type PFN_vkCmdClearDepthStencilImage = fn (command_buffer CommandBuffer, image Image, image_layout ImageLayout, p_depth_stencil &ClearDepthStencilValue, range_count u32, p_ranges &ImageSubresourceRange)

@[inline]
pub fn cmd_clear_depth_stencil_image(command_buffer CommandBuffer,
	image Image,
	image_layout ImageLayout,
	p_depth_stencil &ClearDepthStencilValue,
	range_count u32,
	p_ranges &ImageSubresourceRange) {
	C.vkCmdClearDepthStencilImage(command_buffer, image, image_layout, p_depth_stencil,
		range_count, p_ranges)
}

@[keep_args_alive]
fn C.vkCmdClearAttachments(command_buffer CommandBuffer, attachment_count u32, p_attachments &ClearAttachment, rect_count u32, p_rects &ClearRect)

pub type PFN_vkCmdClearAttachments = fn (command_buffer CommandBuffer, attachment_count u32, p_attachments &ClearAttachment, rect_count u32, p_rects &ClearRect)

@[inline]
pub fn cmd_clear_attachments(command_buffer CommandBuffer,
	attachment_count u32,
	p_attachments &ClearAttachment,
	rect_count u32,
	p_rects &ClearRect) {
	C.vkCmdClearAttachments(command_buffer, attachment_count, p_attachments, rect_count,
		p_rects)
}

@[keep_args_alive]
fn C.vkCmdResolveImage(command_buffer CommandBuffer, src_image Image, src_image_layout ImageLayout, dst_image Image, dst_image_layout ImageLayout, region_count u32, p_regions &ImageResolve)

pub type PFN_vkCmdResolveImage = fn (command_buffer CommandBuffer, src_image Image, src_image_layout ImageLayout, dst_image Image, dst_image_layout ImageLayout, region_count u32, p_regions &ImageResolve)

@[inline]
pub fn cmd_resolve_image(command_buffer CommandBuffer,
	src_image Image,
	src_image_layout ImageLayout,
	dst_image Image,
	dst_image_layout ImageLayout,
	region_count u32,
	p_regions &ImageResolve) {
	C.vkCmdResolveImage(command_buffer, src_image, src_image_layout, dst_image, dst_image_layout,
		region_count, p_regions)
}

@[keep_args_alive]
fn C.vkCmdBeginRenderPass(command_buffer CommandBuffer, p_render_pass_begin &RenderPassBeginInfo, contents SubpassContents)

pub type PFN_vkCmdBeginRenderPass = fn (command_buffer CommandBuffer, p_render_pass_begin &RenderPassBeginInfo, contents SubpassContents)

@[inline]
pub fn cmd_begin_render_pass(command_buffer CommandBuffer,
	p_render_pass_begin &RenderPassBeginInfo,
	contents SubpassContents) {
	C.vkCmdBeginRenderPass(command_buffer, p_render_pass_begin, contents)
}

@[keep_args_alive]
fn C.vkCmdNextSubpass(command_buffer CommandBuffer, contents SubpassContents)

pub type PFN_vkCmdNextSubpass = fn (command_buffer CommandBuffer, contents SubpassContents)

@[inline]
pub fn cmd_next_subpass(command_buffer CommandBuffer,
	contents SubpassContents) {
	C.vkCmdNextSubpass(command_buffer, contents)
}

@[keep_args_alive]
fn C.vkCmdEndRenderPass(command_buffer CommandBuffer)

pub type PFN_vkCmdEndRenderPass = fn (command_buffer CommandBuffer)

@[inline]
pub fn cmd_end_render_pass(command_buffer CommandBuffer) {
	C.vkCmdEndRenderPass(command_buffer)
}

pub const api_version_1_1 = make_api_version(0, 1, 1, 0) // patch version should always be set to 0
// Pointer to VkDescriptorUpdateTemplate_T
pub type DescriptorUpdateTemplate = voidptr

// Pointer to VkSamplerYcbcrConversion_T
pub type SamplerYcbcrConversion = voidptr

pub const max_device_group_size = u32(32)
pub const luid_size = u32(8)
pub const queue_family_external = ~u32(1)

pub enum DescriptorUpdateTemplateType as u32 {
	descriptor_set   = 0
	push_descriptors = 1
	max_enum         = max_int
}

pub enum SamplerYcbcrModelConversion as u32 {
	rgb_identity   = 0
	ycbcr_identity = 1
	ycbcr709       = 2
	ycbcr601       = 3
	ycbcr2020      = 4
	max_enum       = max_int
}

pub enum SamplerYcbcrRange as u32 {
	itu_full   = 0
	itu_narrow = 1
	max_enum   = max_int
}

pub enum ChromaLocation as u32 {
	cosited_even = 0
	midpoint     = 1
	max_enum     = max_int
}

pub enum PointClippingBehavior as u32 {
	all_clip_planes       = 0
	user_clip_planes_only = 1
	max_enum              = max_int
}

pub enum TessellationDomainOrigin as u32 {
	upper_left = 0
	lower_left = 1
	max_enum   = max_int
}

pub enum PeerMemoryFeatureFlagBits as u32 {
	copy_src    = u32(0x00000001)
	copy_dst    = u32(0x00000002)
	generic_src = u32(0x00000004)
	generic_dst = u32(0x00000008)
	max_enum    = max_int
}
pub type PeerMemoryFeatureFlags = u32

pub enum MemoryAllocateFlagBits as u32 {
	device_mask                   = u32(0x00000001)
	device_address                = u32(0x00000002)
	device_address_capture_replay = u32(0x00000004)
	zero_initialize_bit_ext       = u32(0x00000008)
	max_enum                      = max_int
}
pub type MemoryAllocateFlags = u32
pub type CommandPoolTrimFlags = u32

pub enum ExternalMemoryHandleTypeFlagBits as u32 {
	opaque_fd                           = u32(0x00000001)
	opaque_win32                        = u32(0x00000002)
	opaque_win32_kmt                    = u32(0x00000004)
	d3d11_texture                       = u32(0x00000008)
	d3d11_texture_kmt                   = u32(0x00000010)
	d3d12_heap                          = u32(0x00000020)
	d3d12_resource                      = u32(0x00000040)
	dma_buf_bit_ext                     = u32(0x00000200)
	android_hardware_buffer_bit_android = u32(0x00000400)
	host_allocation_bit_ext             = u32(0x00000080)
	host_mapped_foreign_memory_bit_ext  = u32(0x00000100)
	zircon_vmo_bit_fuchsia              = u32(0x00000800)
	rdma_address_bit_nv                 = u32(0x00001000)
	screen_buffer_bit_qnx               = u32(0x00004000)
	mtlbuffer_bit_ext                   = u32(0x00010000)
	mtltexture_bit_ext                  = u32(0x00020000)
	mtlheap_bit_ext                     = u32(0x00040000)
	max_enum                            = max_int
}
pub type ExternalMemoryHandleTypeFlags = u32

pub enum ExternalMemoryFeatureFlagBits as u32 {
	dedicated_only = u32(0x00000001)
	exportable     = u32(0x00000002)
	importable     = u32(0x00000004)
	max_enum       = max_int
}
pub type ExternalMemoryFeatureFlags = u32

pub enum ExternalFenceHandleTypeFlagBits as u32 {
	opaque_fd        = u32(0x00000001)
	opaque_win32     = u32(0x00000002)
	opaque_win32_kmt = u32(0x00000004)
	sync_fd          = u32(0x00000008)
	max_enum         = max_int
}
pub type ExternalFenceHandleTypeFlags = u32

pub enum ExternalFenceFeatureFlagBits as u32 {
	exportable = u32(0x00000001)
	importable = u32(0x00000002)
	max_enum   = max_int
}
pub type ExternalFenceFeatureFlags = u32

pub enum FenceImportFlagBits as u32 {
	temporary = u32(0x00000001)
	max_enum  = max_int
}
pub type FenceImportFlags = u32

pub enum SemaphoreImportFlagBits as u32 {
	temporary = u32(0x00000001)
	max_enum  = max_int
}
pub type SemaphoreImportFlags = u32

pub enum ExternalSemaphoreHandleTypeFlagBits as u32 {
	opaque_fd                = u32(0x00000001)
	opaque_win32             = u32(0x00000002)
	opaque_win32_kmt         = u32(0x00000004)
	d3d12_fence              = u32(0x00000008)
	sync_fd                  = u32(0x00000010)
	zircon_event_bit_fuchsia = u32(0x00000080)
	max_enum                 = max_int
}
pub type ExternalSemaphoreHandleTypeFlags = u32

pub enum ExternalSemaphoreFeatureFlagBits as u32 {
	exportable = u32(0x00000001)
	importable = u32(0x00000002)
	max_enum   = max_int
}
pub type ExternalSemaphoreFeatureFlags = u32

pub enum SubgroupFeatureFlagBits as u32 {
	basic              = u32(0x00000001)
	vote               = u32(0x00000002)
	arithmetic         = u32(0x00000004)
	ballot             = u32(0x00000008)
	shuffle            = u32(0x00000010)
	shuffle_relative   = u32(0x00000020)
	clustered          = u32(0x00000040)
	quad               = u32(0x00000080)
	rotate             = u32(0x00000200)
	rotate_clustered   = u32(0x00000400)
	partitioned_bit_nv = u32(0x00000100)
	max_enum           = max_int
}
pub type SubgroupFeatureFlags = u32
pub type DescriptorUpdateTemplateCreateFlags = u32
pub type BindBufferMemoryInfo = C.VkBindBufferMemoryInfo

@[typedef]
pub struct C.VkBindBufferMemoryInfo {
pub mut:
	sType        StructureType = StructureType.bind_buffer_memory_info
	pNext        voidptr       = unsafe { nil }
	buffer       Buffer
	memory       DeviceMemory
	memoryOffset DeviceSize
}

pub type BindImageMemoryInfo = C.VkBindImageMemoryInfo

@[typedef]
pub struct C.VkBindImageMemoryInfo {
pub mut:
	sType        StructureType = StructureType.bind_image_memory_info
	pNext        voidptr       = unsafe { nil }
	image        Image
	memory       DeviceMemory
	memoryOffset DeviceSize
}

// MemoryDedicatedRequirements extends VkMemoryRequirements2
pub type MemoryDedicatedRequirements = C.VkMemoryDedicatedRequirements

@[typedef]
pub struct C.VkMemoryDedicatedRequirements {
pub mut:
	sType                       StructureType = StructureType.memory_dedicated_requirements
	pNext                       voidptr       = unsafe { nil }
	prefersDedicatedAllocation  Bool32
	requiresDedicatedAllocation Bool32
}

// MemoryDedicatedAllocateInfo extends VkMemoryAllocateInfo
pub type MemoryDedicatedAllocateInfo = C.VkMemoryDedicatedAllocateInfo

@[typedef]
pub struct C.VkMemoryDedicatedAllocateInfo {
pub mut:
	sType  StructureType = StructureType.memory_dedicated_allocate_info
	pNext  voidptr       = unsafe { nil }
	image  Image
	buffer Buffer
}

// MemoryAllocateFlagsInfo extends VkMemoryAllocateInfo
pub type MemoryAllocateFlagsInfo = C.VkMemoryAllocateFlagsInfo

@[typedef]
pub struct C.VkMemoryAllocateFlagsInfo {
pub mut:
	sType      StructureType = StructureType.memory_allocate_flags_info
	pNext      voidptr       = unsafe { nil }
	flags      MemoryAllocateFlags
	deviceMask u32
}

// DeviceGroupCommandBufferBeginInfo extends VkCommandBufferBeginInfo
pub type DeviceGroupCommandBufferBeginInfo = C.VkDeviceGroupCommandBufferBeginInfo

@[typedef]
pub struct C.VkDeviceGroupCommandBufferBeginInfo {
pub mut:
	sType      StructureType = StructureType.device_group_command_buffer_begin_info
	pNext      voidptr       = unsafe { nil }
	deviceMask u32
}

// DeviceGroupSubmitInfo extends VkSubmitInfo
pub type DeviceGroupSubmitInfo = C.VkDeviceGroupSubmitInfo

@[typedef]
pub struct C.VkDeviceGroupSubmitInfo {
pub mut:
	sType                         StructureType = StructureType.device_group_submit_info
	pNext                         voidptr       = unsafe { nil }
	waitSemaphoreCount            u32
	pWaitSemaphoreDeviceIndices   &u32
	commandBufferCount            u32
	pCommandBufferDeviceMasks     &u32
	signalSemaphoreCount          u32
	pSignalSemaphoreDeviceIndices &u32
}

// DeviceGroupBindSparseInfo extends VkBindSparseInfo
pub type DeviceGroupBindSparseInfo = C.VkDeviceGroupBindSparseInfo

@[typedef]
pub struct C.VkDeviceGroupBindSparseInfo {
pub mut:
	sType               StructureType = StructureType.device_group_bind_sparse_info
	pNext               voidptr       = unsafe { nil }
	resourceDeviceIndex u32
	memoryDeviceIndex   u32
}

// BindBufferMemoryDeviceGroupInfo extends VkBindBufferMemoryInfo
pub type BindBufferMemoryDeviceGroupInfo = C.VkBindBufferMemoryDeviceGroupInfo

@[typedef]
pub struct C.VkBindBufferMemoryDeviceGroupInfo {
pub mut:
	sType            StructureType = StructureType.bind_buffer_memory_device_group_info
	pNext            voidptr       = unsafe { nil }
	deviceIndexCount u32
	pDeviceIndices   &u32
}

// BindImageMemoryDeviceGroupInfo extends VkBindImageMemoryInfo
pub type BindImageMemoryDeviceGroupInfo = C.VkBindImageMemoryDeviceGroupInfo

@[typedef]
pub struct C.VkBindImageMemoryDeviceGroupInfo {
pub mut:
	sType                        StructureType = StructureType.bind_image_memory_device_group_info
	pNext                        voidptr       = unsafe { nil }
	deviceIndexCount             u32
	pDeviceIndices               &u32
	splitInstanceBindRegionCount u32
	pSplitInstanceBindRegions    &Rect2D
}

pub type PhysicalDeviceGroupProperties = C.VkPhysicalDeviceGroupProperties

@[typedef]
pub struct C.VkPhysicalDeviceGroupProperties {
pub mut:
	sType               StructureType = StructureType.physical_device_group_properties
	pNext               voidptr       = unsafe { nil }
	physicalDeviceCount u32
	physicalDevices     [max_device_group_size]PhysicalDevice
	subsetAllocation    Bool32
}

// DeviceGroupDeviceCreateInfo extends VkDeviceCreateInfo
pub type DeviceGroupDeviceCreateInfo = C.VkDeviceGroupDeviceCreateInfo

@[typedef]
pub struct C.VkDeviceGroupDeviceCreateInfo {
pub mut:
	sType               StructureType = StructureType.device_group_device_create_info
	pNext               voidptr       = unsafe { nil }
	physicalDeviceCount u32
	pPhysicalDevices    &PhysicalDevice
}

pub type BufferMemoryRequirementsInfo2 = C.VkBufferMemoryRequirementsInfo2

@[typedef]
pub struct C.VkBufferMemoryRequirementsInfo2 {
pub mut:
	sType  StructureType = StructureType.buffer_memory_requirements_info2
	pNext  voidptr       = unsafe { nil }
	buffer Buffer
}

pub type ImageMemoryRequirementsInfo2 = C.VkImageMemoryRequirementsInfo2

@[typedef]
pub struct C.VkImageMemoryRequirementsInfo2 {
pub mut:
	sType StructureType = StructureType.image_memory_requirements_info2
	pNext voidptr       = unsafe { nil }
	image Image
}

pub type ImageSparseMemoryRequirementsInfo2 = C.VkImageSparseMemoryRequirementsInfo2

@[typedef]
pub struct C.VkImageSparseMemoryRequirementsInfo2 {
pub mut:
	sType StructureType = StructureType.image_sparse_memory_requirements_info2
	pNext voidptr       = unsafe { nil }
	image Image
}

pub type MemoryRequirements2 = C.VkMemoryRequirements2

@[typedef]
pub struct C.VkMemoryRequirements2 {
pub mut:
	sType              StructureType = StructureType.memory_requirements2
	pNext              voidptr       = unsafe { nil }
	memoryRequirements MemoryRequirements
}

pub type SparseImageMemoryRequirements2 = C.VkSparseImageMemoryRequirements2

@[typedef]
pub struct C.VkSparseImageMemoryRequirements2 {
pub mut:
	sType              StructureType = StructureType.sparse_image_memory_requirements2
	pNext              voidptr       = unsafe { nil }
	memoryRequirements SparseImageMemoryRequirements
}

// PhysicalDeviceFeatures2 extends VkDeviceCreateInfo
pub type PhysicalDeviceFeatures2 = C.VkPhysicalDeviceFeatures2

@[typedef]
pub struct C.VkPhysicalDeviceFeatures2 {
pub mut:
	sType    StructureType = StructureType.physical_device_features2
	pNext    voidptr       = unsafe { nil }
	features PhysicalDeviceFeatures
}

pub type PhysicalDeviceProperties2 = C.VkPhysicalDeviceProperties2

@[typedef]
pub struct C.VkPhysicalDeviceProperties2 {
pub mut:
	sType      StructureType = StructureType.physical_device_properties2
	pNext      voidptr       = unsafe { nil }
	properties PhysicalDeviceProperties
}

pub type FormatProperties2 = C.VkFormatProperties2

@[typedef]
pub struct C.VkFormatProperties2 {
pub mut:
	sType            StructureType = StructureType.format_properties2
	pNext            voidptr       = unsafe { nil }
	formatProperties FormatProperties
}

pub type ImageFormatProperties2 = C.VkImageFormatProperties2

@[typedef]
pub struct C.VkImageFormatProperties2 {
pub mut:
	sType                 StructureType = StructureType.image_format_properties2
	pNext                 voidptr       = unsafe { nil }
	imageFormatProperties ImageFormatProperties
}

pub type PhysicalDeviceImageFormatInfo2 = C.VkPhysicalDeviceImageFormatInfo2

@[typedef]
pub struct C.VkPhysicalDeviceImageFormatInfo2 {
pub mut:
	sType  StructureType = StructureType.physical_device_image_format_info2
	pNext  voidptr       = unsafe { nil }
	format Format
	type   ImageType
	tiling ImageTiling
	usage  ImageUsageFlags
	flags  ImageCreateFlags
}

pub type QueueFamilyProperties2 = C.VkQueueFamilyProperties2

@[typedef]
pub struct C.VkQueueFamilyProperties2 {
pub mut:
	sType                 StructureType = StructureType.queue_family_properties2
	pNext                 voidptr       = unsafe { nil }
	queueFamilyProperties QueueFamilyProperties
}

pub type PhysicalDeviceMemoryProperties2 = C.VkPhysicalDeviceMemoryProperties2

@[typedef]
pub struct C.VkPhysicalDeviceMemoryProperties2 {
pub mut:
	sType            StructureType = StructureType.physical_device_memory_properties2
	pNext            voidptr       = unsafe { nil }
	memoryProperties PhysicalDeviceMemoryProperties
}

pub type SparseImageFormatProperties2 = C.VkSparseImageFormatProperties2

@[typedef]
pub struct C.VkSparseImageFormatProperties2 {
pub mut:
	sType      StructureType = StructureType.sparse_image_format_properties2
	pNext      voidptr       = unsafe { nil }
	properties SparseImageFormatProperties
}

pub type PhysicalDeviceSparseImageFormatInfo2 = C.VkPhysicalDeviceSparseImageFormatInfo2

@[typedef]
pub struct C.VkPhysicalDeviceSparseImageFormatInfo2 {
pub mut:
	sType   StructureType = StructureType.physical_device_sparse_image_format_info2
	pNext   voidptr       = unsafe { nil }
	format  Format
	type    ImageType
	samples SampleCountFlagBits
	usage   ImageUsageFlags
	tiling  ImageTiling
}

// ImageViewUsageCreateInfo extends VkImageViewCreateInfo
pub type ImageViewUsageCreateInfo = C.VkImageViewUsageCreateInfo

@[typedef]
pub struct C.VkImageViewUsageCreateInfo {
pub mut:
	sType StructureType = StructureType.image_view_usage_create_info
	pNext voidptr       = unsafe { nil }
	usage ImageUsageFlags
}

// PhysicalDeviceProtectedMemoryFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceProtectedMemoryFeatures = C.VkPhysicalDeviceProtectedMemoryFeatures

@[typedef]
pub struct C.VkPhysicalDeviceProtectedMemoryFeatures {
pub mut:
	sType           StructureType = StructureType.physical_device_protected_memory_features
	pNext           voidptr       = unsafe { nil }
	protectedMemory Bool32
}

// PhysicalDeviceProtectedMemoryProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceProtectedMemoryProperties = C.VkPhysicalDeviceProtectedMemoryProperties

@[typedef]
pub struct C.VkPhysicalDeviceProtectedMemoryProperties {
pub mut:
	sType            StructureType = StructureType.physical_device_protected_memory_properties
	pNext            voidptr       = unsafe { nil }
	protectedNoFault Bool32
}

pub type DeviceQueueInfo2 = C.VkDeviceQueueInfo2

@[typedef]
pub struct C.VkDeviceQueueInfo2 {
pub mut:
	sType            StructureType = StructureType.device_queue_info2
	pNext            voidptr       = unsafe { nil }
	flags            DeviceQueueCreateFlags
	queueFamilyIndex u32
	queueIndex       u32
}

// ProtectedSubmitInfo extends VkSubmitInfo
pub type ProtectedSubmitInfo = C.VkProtectedSubmitInfo

@[typedef]
pub struct C.VkProtectedSubmitInfo {
pub mut:
	sType           StructureType = StructureType.protected_submit_info
	pNext           voidptr       = unsafe { nil }
	protectedSubmit Bool32
}

// BindImagePlaneMemoryInfo extends VkBindImageMemoryInfo
pub type BindImagePlaneMemoryInfo = C.VkBindImagePlaneMemoryInfo

@[typedef]
pub struct C.VkBindImagePlaneMemoryInfo {
pub mut:
	sType       StructureType = StructureType.bind_image_plane_memory_info
	pNext       voidptr       = unsafe { nil }
	planeAspect ImageAspectFlagBits
}

// ImagePlaneMemoryRequirementsInfo extends VkImageMemoryRequirementsInfo2
pub type ImagePlaneMemoryRequirementsInfo = C.VkImagePlaneMemoryRequirementsInfo

@[typedef]
pub struct C.VkImagePlaneMemoryRequirementsInfo {
pub mut:
	sType       StructureType = StructureType.image_plane_memory_requirements_info
	pNext       voidptr       = unsafe { nil }
	planeAspect ImageAspectFlagBits
}

pub type ExternalMemoryProperties = C.VkExternalMemoryProperties

@[typedef]
pub struct C.VkExternalMemoryProperties {
pub mut:
	externalMemoryFeatures        ExternalMemoryFeatureFlags
	exportFromImportedHandleTypes ExternalMemoryHandleTypeFlags
	compatibleHandleTypes         ExternalMemoryHandleTypeFlags
}

// PhysicalDeviceExternalImageFormatInfo extends VkPhysicalDeviceImageFormatInfo2
pub type PhysicalDeviceExternalImageFormatInfo = C.VkPhysicalDeviceExternalImageFormatInfo

@[typedef]
pub struct C.VkPhysicalDeviceExternalImageFormatInfo {
pub mut:
	sType      StructureType = StructureType.physical_device_external_image_format_info
	pNext      voidptr       = unsafe { nil }
	handleType ExternalMemoryHandleTypeFlagBits
}

// ExternalImageFormatProperties extends VkImageFormatProperties2
pub type ExternalImageFormatProperties = C.VkExternalImageFormatProperties

@[typedef]
pub struct C.VkExternalImageFormatProperties {
pub mut:
	sType                    StructureType = StructureType.external_image_format_properties
	pNext                    voidptr       = unsafe { nil }
	externalMemoryProperties ExternalMemoryProperties
}

pub type PhysicalDeviceExternalBufferInfo = C.VkPhysicalDeviceExternalBufferInfo

@[typedef]
pub struct C.VkPhysicalDeviceExternalBufferInfo {
pub mut:
	sType      StructureType = StructureType.physical_device_external_buffer_info
	pNext      voidptr       = unsafe { nil }
	flags      BufferCreateFlags
	usage      BufferUsageFlags
	handleType ExternalMemoryHandleTypeFlagBits
}

pub type ExternalBufferProperties = C.VkExternalBufferProperties

@[typedef]
pub struct C.VkExternalBufferProperties {
pub mut:
	sType                    StructureType = StructureType.external_buffer_properties
	pNext                    voidptr       = unsafe { nil }
	externalMemoryProperties ExternalMemoryProperties
}

// PhysicalDeviceIDProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceIDProperties = C.VkPhysicalDeviceIDProperties

@[typedef]
pub struct C.VkPhysicalDeviceIDProperties {
pub mut:
	sType           StructureType = StructureType.physical_device_id_properties
	pNext           voidptr       = unsafe { nil }
	deviceUUID      [uuid_size]u8
	driverUUID      [uuid_size]u8
	deviceLUID      [luid_size]u8
	deviceNodeMask  u32
	deviceLUIDValid Bool32
}

// ExternalMemoryImageCreateInfo extends VkImageCreateInfo
pub type ExternalMemoryImageCreateInfo = C.VkExternalMemoryImageCreateInfo

@[typedef]
pub struct C.VkExternalMemoryImageCreateInfo {
pub mut:
	sType       StructureType = StructureType.external_memory_image_create_info
	pNext       voidptr       = unsafe { nil }
	handleTypes ExternalMemoryHandleTypeFlags
}

// ExternalMemoryBufferCreateInfo extends VkBufferCreateInfo
pub type ExternalMemoryBufferCreateInfo = C.VkExternalMemoryBufferCreateInfo

@[typedef]
pub struct C.VkExternalMemoryBufferCreateInfo {
pub mut:
	sType       StructureType = StructureType.external_memory_buffer_create_info
	pNext       voidptr       = unsafe { nil }
	handleTypes ExternalMemoryHandleTypeFlags
}

// ExportMemoryAllocateInfo extends VkMemoryAllocateInfo
pub type ExportMemoryAllocateInfo = C.VkExportMemoryAllocateInfo

@[typedef]
pub struct C.VkExportMemoryAllocateInfo {
pub mut:
	sType       StructureType = StructureType.export_memory_allocate_info
	pNext       voidptr       = unsafe { nil }
	handleTypes ExternalMemoryHandleTypeFlags
}

pub type PhysicalDeviceExternalFenceInfo = C.VkPhysicalDeviceExternalFenceInfo

@[typedef]
pub struct C.VkPhysicalDeviceExternalFenceInfo {
pub mut:
	sType      StructureType = StructureType.physical_device_external_fence_info
	pNext      voidptr       = unsafe { nil }
	handleType ExternalFenceHandleTypeFlagBits
}

pub type ExternalFenceProperties = C.VkExternalFenceProperties

@[typedef]
pub struct C.VkExternalFenceProperties {
pub mut:
	sType                         StructureType = StructureType.external_fence_properties
	pNext                         voidptr       = unsafe { nil }
	exportFromImportedHandleTypes ExternalFenceHandleTypeFlags
	compatibleHandleTypes         ExternalFenceHandleTypeFlags
	externalFenceFeatures         ExternalFenceFeatureFlags
}

// ExportFenceCreateInfo extends VkFenceCreateInfo
pub type ExportFenceCreateInfo = C.VkExportFenceCreateInfo

@[typedef]
pub struct C.VkExportFenceCreateInfo {
pub mut:
	sType       StructureType = StructureType.export_fence_create_info
	pNext       voidptr       = unsafe { nil }
	handleTypes ExternalFenceHandleTypeFlags
}

// ExportSemaphoreCreateInfo extends VkSemaphoreCreateInfo
pub type ExportSemaphoreCreateInfo = C.VkExportSemaphoreCreateInfo

@[typedef]
pub struct C.VkExportSemaphoreCreateInfo {
pub mut:
	sType       StructureType = StructureType.export_semaphore_create_info
	pNext       voidptr       = unsafe { nil }
	handleTypes ExternalSemaphoreHandleTypeFlags
}

pub type PhysicalDeviceExternalSemaphoreInfo = C.VkPhysicalDeviceExternalSemaphoreInfo

@[typedef]
pub struct C.VkPhysicalDeviceExternalSemaphoreInfo {
pub mut:
	sType      StructureType = StructureType.physical_device_external_semaphore_info
	pNext      voidptr       = unsafe { nil }
	handleType ExternalSemaphoreHandleTypeFlagBits
}

pub type ExternalSemaphoreProperties = C.VkExternalSemaphoreProperties

@[typedef]
pub struct C.VkExternalSemaphoreProperties {
pub mut:
	sType                         StructureType = StructureType.external_semaphore_properties
	pNext                         voidptr       = unsafe { nil }
	exportFromImportedHandleTypes ExternalSemaphoreHandleTypeFlags
	compatibleHandleTypes         ExternalSemaphoreHandleTypeFlags
	externalSemaphoreFeatures     ExternalSemaphoreFeatureFlags
}

// PhysicalDeviceSubgroupProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceSubgroupProperties = C.VkPhysicalDeviceSubgroupProperties

@[typedef]
pub struct C.VkPhysicalDeviceSubgroupProperties {
pub mut:
	sType                     StructureType = StructureType.physical_device_subgroup_properties
	pNext                     voidptr       = unsafe { nil }
	subgroupSize              u32
	supportedStages           ShaderStageFlags
	supportedOperations       SubgroupFeatureFlags
	quadOperationsInAllStages Bool32
}

// PhysicalDevice16BitStorageFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevice16BitStorageFeatures = C.VkPhysicalDevice16BitStorageFeatures

@[typedef]
pub struct C.VkPhysicalDevice16BitStorageFeatures {
pub mut:
	sType                              StructureType = StructureType.physical_device16bit_storage_features
	pNext                              voidptr       = unsafe { nil }
	storageBuffer16BitAccess           Bool32
	uniformAndStorageBuffer16BitAccess Bool32
	storagePushConstant16              Bool32
	storageInputOutput16               Bool32
}

// PhysicalDeviceVariablePointersFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVariablePointersFeatures = C.VkPhysicalDeviceVariablePointersFeatures

@[typedef]
pub struct C.VkPhysicalDeviceVariablePointersFeatures {
pub mut:
	sType                         StructureType = StructureType.physical_device_variable_pointers_features
	pNext                         voidptr       = unsafe { nil }
	variablePointersStorageBuffer Bool32
	variablePointers              Bool32
}

pub type PhysicalDeviceVariablePointerFeatures = C.VkPhysicalDeviceVariablePointersFeatures

pub type DescriptorUpdateTemplateEntry = C.VkDescriptorUpdateTemplateEntry

@[typedef]
pub struct C.VkDescriptorUpdateTemplateEntry {
pub mut:
	dstBinding      u32
	dstArrayElement u32
	descriptorCount u32
	descriptorType  DescriptorType
	offset          usize
	stride          usize
}

pub type DescriptorUpdateTemplateCreateInfo = C.VkDescriptorUpdateTemplateCreateInfo

@[typedef]
pub struct C.VkDescriptorUpdateTemplateCreateInfo {
pub mut:
	sType                      StructureType = StructureType.descriptor_update_template_create_info
	pNext                      voidptr       = unsafe { nil }
	flags                      DescriptorUpdateTemplateCreateFlags
	descriptorUpdateEntryCount u32
	pDescriptorUpdateEntries   &DescriptorUpdateTemplateEntry
	templateType               DescriptorUpdateTemplateType
	descriptorSetLayout        DescriptorSetLayout
	pipelineBindPoint          PipelineBindPoint
	pipelineLayout             PipelineLayout
	set                        u32
}

// PhysicalDeviceMaintenance3Properties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMaintenance3Properties = C.VkPhysicalDeviceMaintenance3Properties

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance3Properties {
pub mut:
	sType                   StructureType = StructureType.physical_device_maintenance3_properties
	pNext                   voidptr       = unsafe { nil }
	maxPerSetDescriptors    u32
	maxMemoryAllocationSize DeviceSize
}

pub type DescriptorSetLayoutSupport = C.VkDescriptorSetLayoutSupport

@[typedef]
pub struct C.VkDescriptorSetLayoutSupport {
pub mut:
	sType     StructureType = StructureType.descriptor_set_layout_support
	pNext     voidptr       = unsafe { nil }
	supported Bool32
}

pub type SamplerYcbcrConversionCreateInfo = C.VkSamplerYcbcrConversionCreateInfo

@[typedef]
pub struct C.VkSamplerYcbcrConversionCreateInfo {
pub mut:
	sType                       StructureType = StructureType.sampler_ycbcr_conversion_create_info
	pNext                       voidptr       = unsafe { nil }
	format                      Format
	ycbcrModel                  SamplerYcbcrModelConversion
	ycbcrRange                  SamplerYcbcrRange
	components                  ComponentMapping
	xChromaOffset               ChromaLocation
	yChromaOffset               ChromaLocation
	chromaFilter                Filter
	forceExplicitReconstruction Bool32
}

// SamplerYcbcrConversionInfo extends VkSamplerCreateInfo,VkImageViewCreateInfo
pub type SamplerYcbcrConversionInfo = C.VkSamplerYcbcrConversionInfo

@[typedef]
pub struct C.VkSamplerYcbcrConversionInfo {
pub mut:
	sType      StructureType = StructureType.sampler_ycbcr_conversion_info
	pNext      voidptr       = unsafe { nil }
	conversion SamplerYcbcrConversion
}

// PhysicalDeviceSamplerYcbcrConversionFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceSamplerYcbcrConversionFeatures = C.VkPhysicalDeviceSamplerYcbcrConversionFeatures

@[typedef]
pub struct C.VkPhysicalDeviceSamplerYcbcrConversionFeatures {
pub mut:
	sType                  StructureType = StructureType.physical_device_sampler_ycbcr_conversion_features
	pNext                  voidptr       = unsafe { nil }
	samplerYcbcrConversion Bool32
}

// SamplerYcbcrConversionImageFormatProperties extends VkImageFormatProperties2
pub type SamplerYcbcrConversionImageFormatProperties = C.VkSamplerYcbcrConversionImageFormatProperties

@[typedef]
pub struct C.VkSamplerYcbcrConversionImageFormatProperties {
pub mut:
	sType                               StructureType = StructureType.sampler_ycbcr_conversion_image_format_properties
	pNext                               voidptr       = unsafe { nil }
	combinedImageSamplerDescriptorCount u32
}

// DeviceGroupRenderPassBeginInfo extends VkRenderPassBeginInfo,VkRenderingInfo
pub type DeviceGroupRenderPassBeginInfo = C.VkDeviceGroupRenderPassBeginInfo

@[typedef]
pub struct C.VkDeviceGroupRenderPassBeginInfo {
pub mut:
	sType                 StructureType = StructureType.device_group_render_pass_begin_info
	pNext                 voidptr       = unsafe { nil }
	deviceMask            u32
	deviceRenderAreaCount u32
	pDeviceRenderAreas    &Rect2D
}

// PhysicalDevicePointClippingProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDevicePointClippingProperties = C.VkPhysicalDevicePointClippingProperties

@[typedef]
pub struct C.VkPhysicalDevicePointClippingProperties {
pub mut:
	sType                 StructureType = StructureType.physical_device_point_clipping_properties
	pNext                 voidptr       = unsafe { nil }
	pointClippingBehavior PointClippingBehavior
}

pub type InputAttachmentAspectReference = C.VkInputAttachmentAspectReference

@[typedef]
pub struct C.VkInputAttachmentAspectReference {
pub mut:
	subpass              u32
	inputAttachmentIndex u32
	aspectMask           ImageAspectFlags
}

// RenderPassInputAttachmentAspectCreateInfo extends VkRenderPassCreateInfo
pub type RenderPassInputAttachmentAspectCreateInfo = C.VkRenderPassInputAttachmentAspectCreateInfo

@[typedef]
pub struct C.VkRenderPassInputAttachmentAspectCreateInfo {
pub mut:
	sType                StructureType = StructureType.render_pass_input_attachment_aspect_create_info
	pNext                voidptr       = unsafe { nil }
	aspectReferenceCount u32
	pAspectReferences    &InputAttachmentAspectReference
}

// PipelineTessellationDomainOriginStateCreateInfo extends VkPipelineTessellationStateCreateInfo
pub type PipelineTessellationDomainOriginStateCreateInfo = C.VkPipelineTessellationDomainOriginStateCreateInfo

@[typedef]
pub struct C.VkPipelineTessellationDomainOriginStateCreateInfo {
pub mut:
	sType        StructureType = StructureType.pipeline_tessellation_domain_origin_state_create_info
	pNext        voidptr       = unsafe { nil }
	domainOrigin TessellationDomainOrigin
}

// RenderPassMultiviewCreateInfo extends VkRenderPassCreateInfo
pub type RenderPassMultiviewCreateInfo = C.VkRenderPassMultiviewCreateInfo

@[typedef]
pub struct C.VkRenderPassMultiviewCreateInfo {
pub mut:
	sType                StructureType = StructureType.render_pass_multiview_create_info
	pNext                voidptr       = unsafe { nil }
	subpassCount         u32
	pViewMasks           &u32
	dependencyCount      u32
	pViewOffsets         &i32
	correlationMaskCount u32
	pCorrelationMasks    &u32
}

// PhysicalDeviceMultiviewFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMultiviewFeatures = C.VkPhysicalDeviceMultiviewFeatures

@[typedef]
pub struct C.VkPhysicalDeviceMultiviewFeatures {
pub mut:
	sType                       StructureType = StructureType.physical_device_multiview_features
	pNext                       voidptr       = unsafe { nil }
	multiview                   Bool32
	multiviewGeometryShader     Bool32
	multiviewTessellationShader Bool32
}

// PhysicalDeviceMultiviewProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMultiviewProperties = C.VkPhysicalDeviceMultiviewProperties

@[typedef]
pub struct C.VkPhysicalDeviceMultiviewProperties {
pub mut:
	sType                     StructureType = StructureType.physical_device_multiview_properties
	pNext                     voidptr       = unsafe { nil }
	maxMultiviewViewCount     u32
	maxMultiviewInstanceIndex u32
}

// PhysicalDeviceShaderDrawParametersFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderDrawParametersFeatures = C.VkPhysicalDeviceShaderDrawParametersFeatures

@[typedef]
pub struct C.VkPhysicalDeviceShaderDrawParametersFeatures {
pub mut:
	sType                StructureType = StructureType.physical_device_shader_draw_parameters_features
	pNext                voidptr       = unsafe { nil }
	shaderDrawParameters Bool32
}

pub type PhysicalDeviceShaderDrawParameterFeatures = C.VkPhysicalDeviceShaderDrawParametersFeatures

@[keep_args_alive]
fn C.vkEnumerateInstanceVersion(p_api_version &u32) Result

pub type PFN_vkEnumerateInstanceVersion = fn (p_api_version &u32) Result

@[inline]
pub fn enumerate_instance_version(p_api_version &u32) Result {
	return C.vkEnumerateInstanceVersion(p_api_version)
}

@[keep_args_alive]
fn C.vkBindBufferMemory2(device Device, bind_info_count u32, p_bind_infos &BindBufferMemoryInfo) Result

pub type PFN_vkBindBufferMemory2 = fn (device Device, bind_info_count u32, p_bind_infos &BindBufferMemoryInfo) Result

@[inline]
pub fn bind_buffer_memory2(device Device,
	bind_info_count u32,
	p_bind_infos &BindBufferMemoryInfo) Result {
	return C.vkBindBufferMemory2(device, bind_info_count, p_bind_infos)
}

@[keep_args_alive]
fn C.vkBindImageMemory2(device Device, bind_info_count u32, p_bind_infos &BindImageMemoryInfo) Result

pub type PFN_vkBindImageMemory2 = fn (device Device, bind_info_count u32, p_bind_infos &BindImageMemoryInfo) Result

@[inline]
pub fn bind_image_memory2(device Device,
	bind_info_count u32,
	p_bind_infos &BindImageMemoryInfo) Result {
	return C.vkBindImageMemory2(device, bind_info_count, p_bind_infos)
}

@[keep_args_alive]
fn C.vkGetDeviceGroupPeerMemoryFeatures(device Device, heap_index u32, local_device_index u32, remote_device_index u32, p_peer_memory_features &PeerMemoryFeatureFlags)

pub type PFN_vkGetDeviceGroupPeerMemoryFeatures = fn (device Device, heap_index u32, local_device_index u32, remote_device_index u32, p_peer_memory_features &PeerMemoryFeatureFlags)

@[inline]
pub fn get_device_group_peer_memory_features(device Device,
	heap_index u32,
	local_device_index u32,
	remote_device_index u32,
	p_peer_memory_features &PeerMemoryFeatureFlags) {
	C.vkGetDeviceGroupPeerMemoryFeatures(device, heap_index, local_device_index, remote_device_index,
		p_peer_memory_features)
}

@[keep_args_alive]
fn C.vkCmdSetDeviceMask(command_buffer CommandBuffer, device_mask u32)

pub type PFN_vkCmdSetDeviceMask = fn (command_buffer CommandBuffer, device_mask u32)

@[inline]
pub fn cmd_set_device_mask(command_buffer CommandBuffer,
	device_mask u32) {
	C.vkCmdSetDeviceMask(command_buffer, device_mask)
}

@[keep_args_alive]
fn C.vkEnumeratePhysicalDeviceGroups(instance Instance, p_physical_device_group_count &u32, mut p_physical_device_group_properties PhysicalDeviceGroupProperties) Result

pub type PFN_vkEnumeratePhysicalDeviceGroups = fn (instance Instance, p_physical_device_group_count &u32, mut p_physical_device_group_properties PhysicalDeviceGroupProperties) Result

@[inline]
pub fn enumerate_physical_device_groups(instance Instance,
	p_physical_device_group_count &u32,
	mut p_physical_device_group_properties PhysicalDeviceGroupProperties) Result {
	return C.vkEnumeratePhysicalDeviceGroups(instance, p_physical_device_group_count, mut
		p_physical_device_group_properties)
}

@[keep_args_alive]
fn C.vkGetImageMemoryRequirements2(device Device, p_info &ImageMemoryRequirementsInfo2, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetImageMemoryRequirements2 = fn (device Device, p_info &ImageMemoryRequirementsInfo2, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_image_memory_requirements2(device Device,
	p_info &ImageMemoryRequirementsInfo2,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetImageMemoryRequirements2(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetBufferMemoryRequirements2(device Device, p_info &BufferMemoryRequirementsInfo2, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetBufferMemoryRequirements2 = fn (device Device, p_info &BufferMemoryRequirementsInfo2, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_buffer_memory_requirements2(device Device,
	p_info &BufferMemoryRequirementsInfo2,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetBufferMemoryRequirements2(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetImageSparseMemoryRequirements2(device Device, p_info &ImageSparseMemoryRequirementsInfo2, p_sparse_memory_requirement_count &u32, mut p_sparse_memory_requirements SparseImageMemoryRequirements2)

pub type PFN_vkGetImageSparseMemoryRequirements2 = fn (device Device, p_info &ImageSparseMemoryRequirementsInfo2, p_sparse_memory_requirement_count &u32, mut p_sparse_memory_requirements SparseImageMemoryRequirements2)

@[inline]
pub fn get_image_sparse_memory_requirements2(device Device,
	p_info &ImageSparseMemoryRequirementsInfo2,
	p_sparse_memory_requirement_count &u32,
	mut p_sparse_memory_requirements SparseImageMemoryRequirements2) {
	C.vkGetImageSparseMemoryRequirements2(device, p_info, p_sparse_memory_requirement_count, mut
		p_sparse_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceFeatures2(physical_device PhysicalDevice, mut p_features PhysicalDeviceFeatures2)

pub type PFN_vkGetPhysicalDeviceFeatures2 = fn (physical_device PhysicalDevice, mut p_features PhysicalDeviceFeatures2)

@[inline]
pub fn get_physical_device_features2(physical_device PhysicalDevice,
	mut p_features PhysicalDeviceFeatures2) {
	C.vkGetPhysicalDeviceFeatures2(physical_device, mut p_features)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceProperties2(physical_device PhysicalDevice, mut p_properties PhysicalDeviceProperties2)

pub type PFN_vkGetPhysicalDeviceProperties2 = fn (physical_device PhysicalDevice, mut p_properties PhysicalDeviceProperties2)

@[inline]
pub fn get_physical_device_properties2(physical_device PhysicalDevice,
	mut p_properties PhysicalDeviceProperties2) {
	C.vkGetPhysicalDeviceProperties2(physical_device, mut p_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceFormatProperties2(physical_device PhysicalDevice, format Format, mut p_format_properties FormatProperties2)

pub type PFN_vkGetPhysicalDeviceFormatProperties2 = fn (physical_device PhysicalDevice, format Format, mut p_format_properties FormatProperties2)

@[inline]
pub fn get_physical_device_format_properties2(physical_device PhysicalDevice,
	format Format,
	mut p_format_properties FormatProperties2) {
	C.vkGetPhysicalDeviceFormatProperties2(physical_device, format, mut p_format_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceImageFormatProperties2(physical_device PhysicalDevice, p_image_format_info &PhysicalDeviceImageFormatInfo2, mut p_image_format_properties ImageFormatProperties2) Result

pub type PFN_vkGetPhysicalDeviceImageFormatProperties2 = fn (physical_device PhysicalDevice, p_image_format_info &PhysicalDeviceImageFormatInfo2, mut p_image_format_properties ImageFormatProperties2) Result

@[inline]
pub fn get_physical_device_image_format_properties2(physical_device PhysicalDevice,
	p_image_format_info &PhysicalDeviceImageFormatInfo2,
	mut p_image_format_properties ImageFormatProperties2) Result {
	return C.vkGetPhysicalDeviceImageFormatProperties2(physical_device, p_image_format_info, mut
		p_image_format_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceQueueFamilyProperties2(physical_device PhysicalDevice, p_queue_family_property_count &u32, mut p_queue_family_properties QueueFamilyProperties2)

pub type PFN_vkGetPhysicalDeviceQueueFamilyProperties2 = fn (physical_device PhysicalDevice, p_queue_family_property_count &u32, mut p_queue_family_properties QueueFamilyProperties2)

@[inline]
pub fn get_physical_device_queue_family_properties2(physical_device PhysicalDevice,
	p_queue_family_property_count &u32,
	mut p_queue_family_properties QueueFamilyProperties2) {
	C.vkGetPhysicalDeviceQueueFamilyProperties2(physical_device, p_queue_family_property_count, mut
		p_queue_family_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceMemoryProperties2(physical_device PhysicalDevice, mut p_memory_properties PhysicalDeviceMemoryProperties2)

pub type PFN_vkGetPhysicalDeviceMemoryProperties2 = fn (physical_device PhysicalDevice, mut p_memory_properties PhysicalDeviceMemoryProperties2)

@[inline]
pub fn get_physical_device_memory_properties2(physical_device PhysicalDevice,
	mut p_memory_properties PhysicalDeviceMemoryProperties2) {
	C.vkGetPhysicalDeviceMemoryProperties2(physical_device, mut p_memory_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceSparseImageFormatProperties2(physical_device PhysicalDevice, p_format_info &PhysicalDeviceSparseImageFormatInfo2, p_property_count &u32, mut p_properties SparseImageFormatProperties2)

pub type PFN_vkGetPhysicalDeviceSparseImageFormatProperties2 = fn (physical_device PhysicalDevice, p_format_info &PhysicalDeviceSparseImageFormatInfo2, p_property_count &u32, mut p_properties SparseImageFormatProperties2)

@[inline]
pub fn get_physical_device_sparse_image_format_properties2(physical_device PhysicalDevice,
	p_format_info &PhysicalDeviceSparseImageFormatInfo2,
	p_property_count &u32,
	mut p_properties SparseImageFormatProperties2) {
	C.vkGetPhysicalDeviceSparseImageFormatProperties2(physical_device, p_format_info,
		p_property_count, mut p_properties)
}

@[keep_args_alive]
fn C.vkTrimCommandPool(device Device, command_pool CommandPool, flags CommandPoolTrimFlags)

pub type PFN_vkTrimCommandPool = fn (device Device, command_pool CommandPool, flags CommandPoolTrimFlags)

@[inline]
pub fn trim_command_pool(device Device,
	command_pool CommandPool,
	flags CommandPoolTrimFlags) {
	C.vkTrimCommandPool(device, command_pool, flags)
}

@[keep_args_alive]
fn C.vkGetDeviceQueue2(device Device, p_queue_info &DeviceQueueInfo2, p_queue &Queue)

pub type PFN_vkGetDeviceQueue2 = fn (device Device, p_queue_info &DeviceQueueInfo2, p_queue &Queue)

@[inline]
pub fn get_device_queue2(device Device,
	p_queue_info &DeviceQueueInfo2,
	p_queue &Queue) {
	C.vkGetDeviceQueue2(device, p_queue_info, p_queue)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceExternalBufferProperties(physical_device PhysicalDevice, p_external_buffer_info &PhysicalDeviceExternalBufferInfo, mut p_external_buffer_properties ExternalBufferProperties)

pub type PFN_vkGetPhysicalDeviceExternalBufferProperties = fn (physical_device PhysicalDevice, p_external_buffer_info &PhysicalDeviceExternalBufferInfo, mut p_external_buffer_properties ExternalBufferProperties)

@[inline]
pub fn get_physical_device_external_buffer_properties(physical_device PhysicalDevice,
	p_external_buffer_info &PhysicalDeviceExternalBufferInfo,
	mut p_external_buffer_properties ExternalBufferProperties) {
	C.vkGetPhysicalDeviceExternalBufferProperties(physical_device, p_external_buffer_info, mut
		p_external_buffer_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceExternalFenceProperties(physical_device PhysicalDevice, p_external_fence_info &PhysicalDeviceExternalFenceInfo, mut p_external_fence_properties ExternalFenceProperties)

pub type PFN_vkGetPhysicalDeviceExternalFenceProperties = fn (physical_device PhysicalDevice, p_external_fence_info &PhysicalDeviceExternalFenceInfo, mut p_external_fence_properties ExternalFenceProperties)

@[inline]
pub fn get_physical_device_external_fence_properties(physical_device PhysicalDevice,
	p_external_fence_info &PhysicalDeviceExternalFenceInfo,
	mut p_external_fence_properties ExternalFenceProperties) {
	C.vkGetPhysicalDeviceExternalFenceProperties(physical_device, p_external_fence_info, mut
		p_external_fence_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceExternalSemaphoreProperties(physical_device PhysicalDevice, p_external_semaphore_info &PhysicalDeviceExternalSemaphoreInfo, mut p_external_semaphore_properties ExternalSemaphoreProperties)

pub type PFN_vkGetPhysicalDeviceExternalSemaphoreProperties = fn (physical_device PhysicalDevice, p_external_semaphore_info &PhysicalDeviceExternalSemaphoreInfo, mut p_external_semaphore_properties ExternalSemaphoreProperties)

@[inline]
pub fn get_physical_device_external_semaphore_properties(physical_device PhysicalDevice,
	p_external_semaphore_info &PhysicalDeviceExternalSemaphoreInfo,
	mut p_external_semaphore_properties ExternalSemaphoreProperties) {
	C.vkGetPhysicalDeviceExternalSemaphoreProperties(physical_device, p_external_semaphore_info, mut
		p_external_semaphore_properties)
}

@[keep_args_alive]
fn C.vkCmdDispatchBase(command_buffer CommandBuffer, base_group_x u32, base_group_y u32, base_group_z u32, group_count_x u32, group_count_y u32, group_count_z u32)

pub type PFN_vkCmdDispatchBase = fn (command_buffer CommandBuffer, base_group_x u32, base_group_y u32, base_group_z u32, group_count_x u32, group_count_y u32, group_count_z u32)

@[inline]
pub fn cmd_dispatch_base(command_buffer CommandBuffer,
	base_group_x u32,
	base_group_y u32,
	base_group_z u32,
	group_count_x u32,
	group_count_y u32,
	group_count_z u32) {
	C.vkCmdDispatchBase(command_buffer, base_group_x, base_group_y, base_group_z, group_count_x,
		group_count_y, group_count_z)
}

@[keep_args_alive]
fn C.vkCreateDescriptorUpdateTemplate(device Device, p_create_info &DescriptorUpdateTemplateCreateInfo, p_allocator &AllocationCallbacks, p_descriptor_update_template &DescriptorUpdateTemplate) Result

pub type PFN_vkCreateDescriptorUpdateTemplate = fn (device Device, p_create_info &DescriptorUpdateTemplateCreateInfo, p_allocator &AllocationCallbacks, p_descriptor_update_template &DescriptorUpdateTemplate) Result

@[inline]
pub fn create_descriptor_update_template(device Device,
	p_create_info &DescriptorUpdateTemplateCreateInfo,
	p_allocator &AllocationCallbacks,
	p_descriptor_update_template &DescriptorUpdateTemplate) Result {
	return C.vkCreateDescriptorUpdateTemplate(device, p_create_info, p_allocator, p_descriptor_update_template)
}

@[keep_args_alive]
fn C.vkDestroyDescriptorUpdateTemplate(device Device, descriptor_update_template DescriptorUpdateTemplate, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyDescriptorUpdateTemplate = fn (device Device, descriptor_update_template DescriptorUpdateTemplate, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_descriptor_update_template(device Device,
	descriptor_update_template DescriptorUpdateTemplate,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyDescriptorUpdateTemplate(device, descriptor_update_template, p_allocator)
}

@[keep_args_alive]
fn C.vkUpdateDescriptorSetWithTemplate(device Device, descriptor_set DescriptorSet, descriptor_update_template DescriptorUpdateTemplate, p_data voidptr)

pub type PFN_vkUpdateDescriptorSetWithTemplate = fn (device Device, descriptor_set DescriptorSet, descriptor_update_template DescriptorUpdateTemplate, p_data voidptr)

@[inline]
pub fn update_descriptor_set_with_template(device Device,
	descriptor_set DescriptorSet,
	descriptor_update_template DescriptorUpdateTemplate,
	p_data voidptr) {
	C.vkUpdateDescriptorSetWithTemplate(device, descriptor_set, descriptor_update_template,
		p_data)
}

@[keep_args_alive]
fn C.vkGetDescriptorSetLayoutSupport(device Device, p_create_info &DescriptorSetLayoutCreateInfo, mut p_support DescriptorSetLayoutSupport)

pub type PFN_vkGetDescriptorSetLayoutSupport = fn (device Device, p_create_info &DescriptorSetLayoutCreateInfo, mut p_support DescriptorSetLayoutSupport)

@[inline]
pub fn get_descriptor_set_layout_support(device Device,
	p_create_info &DescriptorSetLayoutCreateInfo,
	mut p_support DescriptorSetLayoutSupport) {
	C.vkGetDescriptorSetLayoutSupport(device, p_create_info, mut p_support)
}

@[keep_args_alive]
fn C.vkCreateSamplerYcbcrConversion(device Device, p_create_info &SamplerYcbcrConversionCreateInfo, p_allocator &AllocationCallbacks, p_ycbcr_conversion &SamplerYcbcrConversion) Result

pub type PFN_vkCreateSamplerYcbcrConversion = fn (device Device, p_create_info &SamplerYcbcrConversionCreateInfo, p_allocator &AllocationCallbacks, p_ycbcr_conversion &SamplerYcbcrConversion) Result

@[inline]
pub fn create_sampler_ycbcr_conversion(device Device,
	p_create_info &SamplerYcbcrConversionCreateInfo,
	p_allocator &AllocationCallbacks,
	p_ycbcr_conversion &SamplerYcbcrConversion) Result {
	return C.vkCreateSamplerYcbcrConversion(device, p_create_info, p_allocator, p_ycbcr_conversion)
}

@[keep_args_alive]
fn C.vkDestroySamplerYcbcrConversion(device Device, ycbcr_conversion SamplerYcbcrConversion, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroySamplerYcbcrConversion = fn (device Device, ycbcr_conversion SamplerYcbcrConversion, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_sampler_ycbcr_conversion(device Device,
	ycbcr_conversion SamplerYcbcrConversion,
	p_allocator &AllocationCallbacks) {
	C.vkDestroySamplerYcbcrConversion(device, ycbcr_conversion, p_allocator)
}

pub const api_version_1_2 = make_api_version(0, 1, 2, 0) // patch version should always be set to 0
pub const max_driver_name_size = u32(256)
pub const max_driver_info_size = u32(256)

pub enum DriverId as u32 {
	amd_proprietary               = 1
	amd_open_source               = 2
	mesa_radv                     = 3
	nvidia_proprietary            = 4
	intel_proprietary_windows     = 5
	intel_open_source_mesa        = 6
	imagination_proprietary       = 7
	qualcomm_proprietary          = 8
	arm_proprietary               = 9
	google_swiftshader            = 10
	ggp_proprietary               = 11
	broadcom_proprietary          = 12
	mesa_llvmpipe                 = 13
	moltenvk                      = 14
	coreavi_proprietary           = 15
	juice_proprietary             = 16
	verisilicon_proprietary       = 17
	mesa_turnip                   = 18
	mesa_v3dv                     = 19
	mesa_panvk                    = 20
	samsung_proprietary           = 21
	mesa_venus                    = 22
	mesa_dozen                    = 23
	mesa_nvk                      = 24
	imagination_open_source_mesa  = 25
	mesa_honeykrisp               = 26
	vulkan_sc_emulation_on_vulkan = 27
	mesa_kosmickrisp              = 28
	max_enum                      = max_int
}

pub enum ShaderFloatControlsIndependence as u32 {
	_32_bit_only = 0
	all          = 1
	none         = 2
	max_enum     = max_int
}

pub enum SemaphoreType as u32 {
	binary   = 0
	timeline = 1
	max_enum = max_int
}

pub enum SamplerReductionMode as u32 {
	weighted_average                 = 0
	min                              = 1
	max                              = 2
	weighted_average_rangeclamp_qcom = 1000521000
	max_enum                         = max_int
}

pub enum ResolveModeFlagBits as u32 {
	none                                   = 0
	sample_zero                            = u32(0x00000001)
	average                                = u32(0x00000002)
	min                                    = u32(0x00000004)
	max                                    = u32(0x00000008)
	external_format_downsample_bit_android = u32(0x00000010)
	max_enum                               = max_int
}
pub type ResolveModeFlags = u32

pub enum SemaphoreWaitFlagBits as u32 {
	any      = u32(0x00000001)
	max_enum = max_int
}
pub type SemaphoreWaitFlags = u32

pub enum DescriptorBindingFlagBits as u32 {
	update_after_bind           = u32(0x00000001)
	update_unused_while_pending = u32(0x00000002)
	partially_bound             = u32(0x00000004)
	variable_descriptor_count   = u32(0x00000008)
	max_enum                    = max_int
}
pub type DescriptorBindingFlags = u32

// PhysicalDeviceVulkan11Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVulkan11Features = C.VkPhysicalDeviceVulkan11Features

@[typedef]
pub struct C.VkPhysicalDeviceVulkan11Features {
pub mut:
	sType                              StructureType = StructureType.physical_device_vulkan1_1_features
	pNext                              voidptr       = unsafe { nil }
	storageBuffer16BitAccess           Bool32
	uniformAndStorageBuffer16BitAccess Bool32
	storagePushConstant16              Bool32
	storageInputOutput16               Bool32
	multiview                          Bool32
	multiviewGeometryShader            Bool32
	multiviewTessellationShader        Bool32
	variablePointersStorageBuffer      Bool32
	variablePointers                   Bool32
	protectedMemory                    Bool32
	samplerYcbcrConversion             Bool32
	shaderDrawParameters               Bool32
}

// PhysicalDeviceVulkan11Properties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceVulkan11Properties = C.VkPhysicalDeviceVulkan11Properties

@[typedef]
pub struct C.VkPhysicalDeviceVulkan11Properties {
pub mut:
	sType                             StructureType = StructureType.physical_device_vulkan1_1_properties
	pNext                             voidptr       = unsafe { nil }
	deviceUUID                        [uuid_size]u8
	driverUUID                        [uuid_size]u8
	deviceLUID                        [luid_size]u8
	deviceNodeMask                    u32
	deviceLUIDValid                   Bool32
	subgroupSize                      u32
	subgroupSupportedStages           ShaderStageFlags
	subgroupSupportedOperations       SubgroupFeatureFlags
	subgroupQuadOperationsInAllStages Bool32
	pointClippingBehavior             PointClippingBehavior
	maxMultiviewViewCount             u32
	maxMultiviewInstanceIndex         u32
	protectedNoFault                  Bool32
	maxPerSetDescriptors              u32
	maxMemoryAllocationSize           DeviceSize
}

// PhysicalDeviceVulkan12Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVulkan12Features = C.VkPhysicalDeviceVulkan12Features

@[typedef]
pub struct C.VkPhysicalDeviceVulkan12Features {
pub mut:
	sType                                              StructureType = StructureType.physical_device_vulkan1_2_features
	pNext                                              voidptr       = unsafe { nil }
	samplerMirrorClampToEdge                           Bool32
	drawIndirectCount                                  Bool32
	storageBuffer8BitAccess                            Bool32
	uniformAndStorageBuffer8BitAccess                  Bool32
	storagePushConstant8                               Bool32
	shaderBufferInt64Atomics                           Bool32
	shaderSharedInt64Atomics                           Bool32
	shaderFloat16                                      Bool32
	shaderInt8                                         Bool32
	descriptorIndexing                                 Bool32
	shaderInputAttachmentArrayDynamicIndexing          Bool32
	shaderUniformTexelBufferArrayDynamicIndexing       Bool32
	shaderStorageTexelBufferArrayDynamicIndexing       Bool32
	shaderUniformBufferArrayNonUniformIndexing         Bool32
	shaderSampledImageArrayNonUniformIndexing          Bool32
	shaderStorageBufferArrayNonUniformIndexing         Bool32
	shaderStorageImageArrayNonUniformIndexing          Bool32
	shaderInputAttachmentArrayNonUniformIndexing       Bool32
	shaderUniformTexelBufferArrayNonUniformIndexing    Bool32
	shaderStorageTexelBufferArrayNonUniformIndexing    Bool32
	descriptorBindingUniformBufferUpdateAfterBind      Bool32
	descriptorBindingSampledImageUpdateAfterBind       Bool32
	descriptorBindingStorageImageUpdateAfterBind       Bool32
	descriptorBindingStorageBufferUpdateAfterBind      Bool32
	descriptorBindingUniformTexelBufferUpdateAfterBind Bool32
	descriptorBindingStorageTexelBufferUpdateAfterBind Bool32
	descriptorBindingUpdateUnusedWhilePending          Bool32
	descriptorBindingPartiallyBound                    Bool32
	descriptorBindingVariableDescriptorCount           Bool32
	runtimeDescriptorArray                             Bool32
	samplerFilterMinmax                                Bool32
	scalarBlockLayout                                  Bool32
	imagelessFramebuffer                               Bool32
	uniformBufferStandardLayout                        Bool32
	shaderSubgroupExtendedTypes                        Bool32
	separateDepthStencilLayouts                        Bool32
	hostQueryReset                                     Bool32
	timelineSemaphore                                  Bool32
	bufferDeviceAddress                                Bool32
	bufferDeviceAddressCaptureReplay                   Bool32
	bufferDeviceAddressMultiDevice                     Bool32
	vulkanMemoryModel                                  Bool32
	vulkanMemoryModelDeviceScope                       Bool32
	vulkanMemoryModelAvailabilityVisibilityChains      Bool32
	shaderOutputViewportIndex                          Bool32
	shaderOutputLayer                                  Bool32
	subgroupBroadcastDynamicId                         Bool32
}

pub type ConformanceVersion = C.VkConformanceVersion

@[typedef]
pub struct C.VkConformanceVersion {
pub mut:
	major    u8
	minor    u8
	subminor u8
	patch    u8
}

// PhysicalDeviceVulkan12Properties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceVulkan12Properties = C.VkPhysicalDeviceVulkan12Properties

@[typedef]
pub struct C.VkPhysicalDeviceVulkan12Properties {
pub mut:
	sType                                                StructureType = StructureType.physical_device_vulkan1_2_properties
	pNext                                                voidptr       = unsafe { nil }
	driverID                                             DriverId
	driverName                                           [max_driver_name_size]char
	driverInfo                                           [max_driver_info_size]char
	conformanceVersion                                   ConformanceVersion
	denormBehaviorIndependence                           ShaderFloatControlsIndependence
	roundingModeIndependence                             ShaderFloatControlsIndependence
	shaderSignedZeroInfNanPreserveFloat16                Bool32
	shaderSignedZeroInfNanPreserveFloat32                Bool32
	shaderSignedZeroInfNanPreserveFloat64                Bool32
	shaderDenormPreserveFloat16                          Bool32
	shaderDenormPreserveFloat32                          Bool32
	shaderDenormPreserveFloat64                          Bool32
	shaderDenormFlushToZeroFloat16                       Bool32
	shaderDenormFlushToZeroFloat32                       Bool32
	shaderDenormFlushToZeroFloat64                       Bool32
	shaderRoundingModeRTEFloat16                         Bool32
	shaderRoundingModeRTEFloat32                         Bool32
	shaderRoundingModeRTEFloat64                         Bool32
	shaderRoundingModeRTZFloat16                         Bool32
	shaderRoundingModeRTZFloat32                         Bool32
	shaderRoundingModeRTZFloat64                         Bool32
	maxUpdateAfterBindDescriptorsInAllPools              u32
	shaderUniformBufferArrayNonUniformIndexingNative     Bool32
	shaderSampledImageArrayNonUniformIndexingNative      Bool32
	shaderStorageBufferArrayNonUniformIndexingNative     Bool32
	shaderStorageImageArrayNonUniformIndexingNative      Bool32
	shaderInputAttachmentArrayNonUniformIndexingNative   Bool32
	robustBufferAccessUpdateAfterBind                    Bool32
	quadDivergentImplicitLod                             Bool32
	maxPerStageDescriptorUpdateAfterBindSamplers         u32
	maxPerStageDescriptorUpdateAfterBindUniformBuffers   u32
	maxPerStageDescriptorUpdateAfterBindStorageBuffers   u32
	maxPerStageDescriptorUpdateAfterBindSampledImages    u32
	maxPerStageDescriptorUpdateAfterBindStorageImages    u32
	maxPerStageDescriptorUpdateAfterBindInputAttachments u32
	maxPerStageUpdateAfterBindResources                  u32
	maxDescriptorSetUpdateAfterBindSamplers              u32
	maxDescriptorSetUpdateAfterBindUniformBuffers        u32
	maxDescriptorSetUpdateAfterBindUniformBuffersDynamic u32
	maxDescriptorSetUpdateAfterBindStorageBuffers        u32
	maxDescriptorSetUpdateAfterBindStorageBuffersDynamic u32
	maxDescriptorSetUpdateAfterBindSampledImages         u32
	maxDescriptorSetUpdateAfterBindStorageImages         u32
	maxDescriptorSetUpdateAfterBindInputAttachments      u32
	supportedDepthResolveModes                           ResolveModeFlags
	supportedStencilResolveModes                         ResolveModeFlags
	independentResolveNone                               Bool32
	independentResolve                                   Bool32
	filterMinmaxSingleComponentFormats                   Bool32
	filterMinmaxImageComponentMapping                    Bool32
	maxTimelineSemaphoreValueDifference                  u64
	framebufferIntegerColorSampleCounts                  SampleCountFlags
}

// ImageFormatListCreateInfo extends VkImageCreateInfo,VkSwapchainCreateInfoKHR,VkPhysicalDeviceImageFormatInfo2
pub type ImageFormatListCreateInfo = C.VkImageFormatListCreateInfo

@[typedef]
pub struct C.VkImageFormatListCreateInfo {
pub mut:
	sType           StructureType = StructureType.image_format_list_create_info
	pNext           voidptr       = unsafe { nil }
	viewFormatCount u32
	pViewFormats    &Format
}

// PhysicalDeviceDriverProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceDriverProperties = C.VkPhysicalDeviceDriverProperties

@[typedef]
pub struct C.VkPhysicalDeviceDriverProperties {
pub mut:
	sType              StructureType = StructureType.physical_device_driver_properties
	pNext              voidptr       = unsafe { nil }
	driverID           DriverId
	driverName         [max_driver_name_size]char
	driverInfo         [max_driver_info_size]char
	conformanceVersion ConformanceVersion
}

// PhysicalDeviceVulkanMemoryModelFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVulkanMemoryModelFeatures = C.VkPhysicalDeviceVulkanMemoryModelFeatures

@[typedef]
pub struct C.VkPhysicalDeviceVulkanMemoryModelFeatures {
pub mut:
	sType                                         StructureType = StructureType.physical_device_vulkan_memory_model_features
	pNext                                         voidptr       = unsafe { nil }
	vulkanMemoryModel                             Bool32
	vulkanMemoryModelDeviceScope                  Bool32
	vulkanMemoryModelAvailabilityVisibilityChains Bool32
}

// PhysicalDeviceHostQueryResetFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceHostQueryResetFeatures = C.VkPhysicalDeviceHostQueryResetFeatures

@[typedef]
pub struct C.VkPhysicalDeviceHostQueryResetFeatures {
pub mut:
	sType          StructureType = StructureType.physical_device_host_query_reset_features
	pNext          voidptr       = unsafe { nil }
	hostQueryReset Bool32
}

// PhysicalDeviceTimelineSemaphoreFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceTimelineSemaphoreFeatures = C.VkPhysicalDeviceTimelineSemaphoreFeatures

@[typedef]
pub struct C.VkPhysicalDeviceTimelineSemaphoreFeatures {
pub mut:
	sType             StructureType = StructureType.physical_device_timeline_semaphore_features
	pNext             voidptr       = unsafe { nil }
	timelineSemaphore Bool32
}

// PhysicalDeviceTimelineSemaphoreProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceTimelineSemaphoreProperties = C.VkPhysicalDeviceTimelineSemaphoreProperties

@[typedef]
pub struct C.VkPhysicalDeviceTimelineSemaphoreProperties {
pub mut:
	sType                               StructureType = StructureType.physical_device_timeline_semaphore_properties
	pNext                               voidptr       = unsafe { nil }
	maxTimelineSemaphoreValueDifference u64
}

// SemaphoreTypeCreateInfo extends VkSemaphoreCreateInfo,VkPhysicalDeviceExternalSemaphoreInfo
pub type SemaphoreTypeCreateInfo = C.VkSemaphoreTypeCreateInfo

@[typedef]
pub struct C.VkSemaphoreTypeCreateInfo {
pub mut:
	sType         StructureType = StructureType.semaphore_type_create_info
	pNext         voidptr       = unsafe { nil }
	semaphoreType SemaphoreType
	initialValue  u64
}

// TimelineSemaphoreSubmitInfo extends VkSubmitInfo,VkBindSparseInfo
pub type TimelineSemaphoreSubmitInfo = C.VkTimelineSemaphoreSubmitInfo

@[typedef]
pub struct C.VkTimelineSemaphoreSubmitInfo {
pub mut:
	sType                     StructureType = StructureType.timeline_semaphore_submit_info
	pNext                     voidptr       = unsafe { nil }
	waitSemaphoreValueCount   u32
	pWaitSemaphoreValues      &u64
	signalSemaphoreValueCount u32
	pSignalSemaphoreValues    &u64
}

pub type SemaphoreWaitInfo = C.VkSemaphoreWaitInfo

@[typedef]
pub struct C.VkSemaphoreWaitInfo {
pub mut:
	sType          StructureType = StructureType.semaphore_wait_info
	pNext          voidptr       = unsafe { nil }
	flags          SemaphoreWaitFlags
	semaphoreCount u32
	pSemaphores    &Semaphore
	pValues        &u64
}

pub type SemaphoreSignalInfo = C.VkSemaphoreSignalInfo

@[typedef]
pub struct C.VkSemaphoreSignalInfo {
pub mut:
	sType     StructureType = StructureType.semaphore_signal_info
	pNext     voidptr       = unsafe { nil }
	semaphore Semaphore
	value     u64
}

// PhysicalDeviceBufferDeviceAddressFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceBufferDeviceAddressFeatures = C.VkPhysicalDeviceBufferDeviceAddressFeatures

@[typedef]
pub struct C.VkPhysicalDeviceBufferDeviceAddressFeatures {
pub mut:
	sType                            StructureType = StructureType.physical_device_buffer_device_address_features
	pNext                            voidptr       = unsafe { nil }
	bufferDeviceAddress              Bool32
	bufferDeviceAddressCaptureReplay Bool32
	bufferDeviceAddressMultiDevice   Bool32
}

pub type BufferDeviceAddressInfo = C.VkBufferDeviceAddressInfo

@[typedef]
pub struct C.VkBufferDeviceAddressInfo {
pub mut:
	sType  StructureType = StructureType.buffer_device_address_info
	pNext  voidptr       = unsafe { nil }
	buffer Buffer
}

// BufferOpaqueCaptureAddressCreateInfo extends VkBufferCreateInfo
pub type BufferOpaqueCaptureAddressCreateInfo = C.VkBufferOpaqueCaptureAddressCreateInfo

@[typedef]
pub struct C.VkBufferOpaqueCaptureAddressCreateInfo {
pub mut:
	sType                StructureType = StructureType.buffer_opaque_capture_address_create_info
	pNext                voidptr       = unsafe { nil }
	opaqueCaptureAddress u64
}

// MemoryOpaqueCaptureAddressAllocateInfo extends VkMemoryAllocateInfo
pub type MemoryOpaqueCaptureAddressAllocateInfo = C.VkMemoryOpaqueCaptureAddressAllocateInfo

@[typedef]
pub struct C.VkMemoryOpaqueCaptureAddressAllocateInfo {
pub mut:
	sType                StructureType = StructureType.memory_opaque_capture_address_allocate_info
	pNext                voidptr       = unsafe { nil }
	opaqueCaptureAddress u64
}

pub type DeviceMemoryOpaqueCaptureAddressInfo = C.VkDeviceMemoryOpaqueCaptureAddressInfo

@[typedef]
pub struct C.VkDeviceMemoryOpaqueCaptureAddressInfo {
pub mut:
	sType  StructureType = StructureType.device_memory_opaque_capture_address_info
	pNext  voidptr       = unsafe { nil }
	memory DeviceMemory
}

// PhysicalDevice8BitStorageFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevice8BitStorageFeatures = C.VkPhysicalDevice8BitStorageFeatures

@[typedef]
pub struct C.VkPhysicalDevice8BitStorageFeatures {
pub mut:
	sType                             StructureType = StructureType.physical_device8bit_storage_features
	pNext                             voidptr       = unsafe { nil }
	storageBuffer8BitAccess           Bool32
	uniformAndStorageBuffer8BitAccess Bool32
	storagePushConstant8              Bool32
}

// PhysicalDeviceShaderAtomicInt64Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderAtomicInt64Features = C.VkPhysicalDeviceShaderAtomicInt64Features

@[typedef]
pub struct C.VkPhysicalDeviceShaderAtomicInt64Features {
pub mut:
	sType                    StructureType = StructureType.physical_device_shader_atomic_int64_features
	pNext                    voidptr       = unsafe { nil }
	shaderBufferInt64Atomics Bool32
	shaderSharedInt64Atomics Bool32
}

// PhysicalDeviceShaderFloat16Int8Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderFloat16Int8Features = C.VkPhysicalDeviceShaderFloat16Int8Features

@[typedef]
pub struct C.VkPhysicalDeviceShaderFloat16Int8Features {
pub mut:
	sType         StructureType = StructureType.physical_device_shader_float16_int8_features
	pNext         voidptr       = unsafe { nil }
	shaderFloat16 Bool32
	shaderInt8    Bool32
}

// PhysicalDeviceFloatControlsProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceFloatControlsProperties = C.VkPhysicalDeviceFloatControlsProperties

@[typedef]
pub struct C.VkPhysicalDeviceFloatControlsProperties {
pub mut:
	sType                                 StructureType = StructureType.physical_device_float_controls_properties
	pNext                                 voidptr       = unsafe { nil }
	denormBehaviorIndependence            ShaderFloatControlsIndependence
	roundingModeIndependence              ShaderFloatControlsIndependence
	shaderSignedZeroInfNanPreserveFloat16 Bool32
	shaderSignedZeroInfNanPreserveFloat32 Bool32
	shaderSignedZeroInfNanPreserveFloat64 Bool32
	shaderDenormPreserveFloat16           Bool32
	shaderDenormPreserveFloat32           Bool32
	shaderDenormPreserveFloat64           Bool32
	shaderDenormFlushToZeroFloat16        Bool32
	shaderDenormFlushToZeroFloat32        Bool32
	shaderDenormFlushToZeroFloat64        Bool32
	shaderRoundingModeRTEFloat16          Bool32
	shaderRoundingModeRTEFloat32          Bool32
	shaderRoundingModeRTEFloat64          Bool32
	shaderRoundingModeRTZFloat16          Bool32
	shaderRoundingModeRTZFloat32          Bool32
	shaderRoundingModeRTZFloat64          Bool32
}

// DescriptorSetLayoutBindingFlagsCreateInfo extends VkDescriptorSetLayoutCreateInfo
pub type DescriptorSetLayoutBindingFlagsCreateInfo = C.VkDescriptorSetLayoutBindingFlagsCreateInfo

@[typedef]
pub struct C.VkDescriptorSetLayoutBindingFlagsCreateInfo {
pub mut:
	sType         StructureType = StructureType.descriptor_set_layout_binding_flags_create_info
	pNext         voidptr       = unsafe { nil }
	bindingCount  u32
	pBindingFlags &DescriptorBindingFlags
}

// PhysicalDeviceDescriptorIndexingFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDescriptorIndexingFeatures = C.VkPhysicalDeviceDescriptorIndexingFeatures

@[typedef]
pub struct C.VkPhysicalDeviceDescriptorIndexingFeatures {
pub mut:
	sType                                              StructureType = StructureType.physical_device_descriptor_indexing_features
	pNext                                              voidptr       = unsafe { nil }
	shaderInputAttachmentArrayDynamicIndexing          Bool32
	shaderUniformTexelBufferArrayDynamicIndexing       Bool32
	shaderStorageTexelBufferArrayDynamicIndexing       Bool32
	shaderUniformBufferArrayNonUniformIndexing         Bool32
	shaderSampledImageArrayNonUniformIndexing          Bool32
	shaderStorageBufferArrayNonUniformIndexing         Bool32
	shaderStorageImageArrayNonUniformIndexing          Bool32
	shaderInputAttachmentArrayNonUniformIndexing       Bool32
	shaderUniformTexelBufferArrayNonUniformIndexing    Bool32
	shaderStorageTexelBufferArrayNonUniformIndexing    Bool32
	descriptorBindingUniformBufferUpdateAfterBind      Bool32
	descriptorBindingSampledImageUpdateAfterBind       Bool32
	descriptorBindingStorageImageUpdateAfterBind       Bool32
	descriptorBindingStorageBufferUpdateAfterBind      Bool32
	descriptorBindingUniformTexelBufferUpdateAfterBind Bool32
	descriptorBindingStorageTexelBufferUpdateAfterBind Bool32
	descriptorBindingUpdateUnusedWhilePending          Bool32
	descriptorBindingPartiallyBound                    Bool32
	descriptorBindingVariableDescriptorCount           Bool32
	runtimeDescriptorArray                             Bool32
}

// PhysicalDeviceDescriptorIndexingProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceDescriptorIndexingProperties = C.VkPhysicalDeviceDescriptorIndexingProperties

@[typedef]
pub struct C.VkPhysicalDeviceDescriptorIndexingProperties {
pub mut:
	sType                                                StructureType = StructureType.physical_device_descriptor_indexing_properties
	pNext                                                voidptr       = unsafe { nil }
	maxUpdateAfterBindDescriptorsInAllPools              u32
	shaderUniformBufferArrayNonUniformIndexingNative     Bool32
	shaderSampledImageArrayNonUniformIndexingNative      Bool32
	shaderStorageBufferArrayNonUniformIndexingNative     Bool32
	shaderStorageImageArrayNonUniformIndexingNative      Bool32
	shaderInputAttachmentArrayNonUniformIndexingNative   Bool32
	robustBufferAccessUpdateAfterBind                    Bool32
	quadDivergentImplicitLod                             Bool32
	maxPerStageDescriptorUpdateAfterBindSamplers         u32
	maxPerStageDescriptorUpdateAfterBindUniformBuffers   u32
	maxPerStageDescriptorUpdateAfterBindStorageBuffers   u32
	maxPerStageDescriptorUpdateAfterBindSampledImages    u32
	maxPerStageDescriptorUpdateAfterBindStorageImages    u32
	maxPerStageDescriptorUpdateAfterBindInputAttachments u32
	maxPerStageUpdateAfterBindResources                  u32
	maxDescriptorSetUpdateAfterBindSamplers              u32
	maxDescriptorSetUpdateAfterBindUniformBuffers        u32
	maxDescriptorSetUpdateAfterBindUniformBuffersDynamic u32
	maxDescriptorSetUpdateAfterBindStorageBuffers        u32
	maxDescriptorSetUpdateAfterBindStorageBuffersDynamic u32
	maxDescriptorSetUpdateAfterBindSampledImages         u32
	maxDescriptorSetUpdateAfterBindStorageImages         u32
	maxDescriptorSetUpdateAfterBindInputAttachments      u32
}

// DescriptorSetVariableDescriptorCountAllocateInfo extends VkDescriptorSetAllocateInfo
pub type DescriptorSetVariableDescriptorCountAllocateInfo = C.VkDescriptorSetVariableDescriptorCountAllocateInfo

@[typedef]
pub struct C.VkDescriptorSetVariableDescriptorCountAllocateInfo {
pub mut:
	sType              StructureType = StructureType.descriptor_set_variable_descriptor_count_allocate_info
	pNext              voidptr       = unsafe { nil }
	descriptorSetCount u32
	pDescriptorCounts  &u32
}

// DescriptorSetVariableDescriptorCountLayoutSupport extends VkDescriptorSetLayoutSupport
pub type DescriptorSetVariableDescriptorCountLayoutSupport = C.VkDescriptorSetVariableDescriptorCountLayoutSupport

@[typedef]
pub struct C.VkDescriptorSetVariableDescriptorCountLayoutSupport {
pub mut:
	sType                      StructureType = StructureType.descriptor_set_variable_descriptor_count_layout_support
	pNext                      voidptr       = unsafe { nil }
	maxVariableDescriptorCount u32
}

// PhysicalDeviceScalarBlockLayoutFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceScalarBlockLayoutFeatures = C.VkPhysicalDeviceScalarBlockLayoutFeatures

@[typedef]
pub struct C.VkPhysicalDeviceScalarBlockLayoutFeatures {
pub mut:
	sType             StructureType = StructureType.physical_device_scalar_block_layout_features
	pNext             voidptr       = unsafe { nil }
	scalarBlockLayout Bool32
}

// SamplerReductionModeCreateInfo extends VkSamplerCreateInfo
pub type SamplerReductionModeCreateInfo = C.VkSamplerReductionModeCreateInfo

@[typedef]
pub struct C.VkSamplerReductionModeCreateInfo {
pub mut:
	sType         StructureType = StructureType.sampler_reduction_mode_create_info
	pNext         voidptr       = unsafe { nil }
	reductionMode SamplerReductionMode
}

// PhysicalDeviceSamplerFilterMinmaxProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceSamplerFilterMinmaxProperties = C.VkPhysicalDeviceSamplerFilterMinmaxProperties

@[typedef]
pub struct C.VkPhysicalDeviceSamplerFilterMinmaxProperties {
pub mut:
	sType                              StructureType = StructureType.physical_device_sampler_filter_minmax_properties
	pNext                              voidptr       = unsafe { nil }
	filterMinmaxSingleComponentFormats Bool32
	filterMinmaxImageComponentMapping  Bool32
}

// PhysicalDeviceUniformBufferStandardLayoutFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceUniformBufferStandardLayoutFeatures = C.VkPhysicalDeviceUniformBufferStandardLayoutFeatures

@[typedef]
pub struct C.VkPhysicalDeviceUniformBufferStandardLayoutFeatures {
pub mut:
	sType                       StructureType = StructureType.physical_device_uniform_buffer_standard_layout_features
	pNext                       voidptr       = unsafe { nil }
	uniformBufferStandardLayout Bool32
}

// PhysicalDeviceShaderSubgroupExtendedTypesFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderSubgroupExtendedTypesFeatures = C.VkPhysicalDeviceShaderSubgroupExtendedTypesFeatures

@[typedef]
pub struct C.VkPhysicalDeviceShaderSubgroupExtendedTypesFeatures {
pub mut:
	sType                       StructureType = StructureType.physical_device_shader_subgroup_extended_types_features
	pNext                       voidptr       = unsafe { nil }
	shaderSubgroupExtendedTypes Bool32
}

pub type AttachmentDescription2 = C.VkAttachmentDescription2

@[typedef]
pub struct C.VkAttachmentDescription2 {
pub mut:
	sType          StructureType = StructureType.attachment_description2
	pNext          voidptr       = unsafe { nil }
	flags          AttachmentDescriptionFlags
	format         Format
	samples        SampleCountFlagBits
	loadOp         AttachmentLoadOp
	storeOp        AttachmentStoreOp
	stencilLoadOp  AttachmentLoadOp
	stencilStoreOp AttachmentStoreOp
	initialLayout  ImageLayout
	finalLayout    ImageLayout
}

pub type AttachmentReference2 = C.VkAttachmentReference2

@[typedef]
pub struct C.VkAttachmentReference2 {
pub mut:
	sType      StructureType = StructureType.attachment_reference2
	pNext      voidptr       = unsafe { nil }
	attachment u32
	layout     ImageLayout
	aspectMask ImageAspectFlags
}

pub type SubpassDescription2 = C.VkSubpassDescription2

@[typedef]
pub struct C.VkSubpassDescription2 {
pub mut:
	sType                   StructureType = StructureType.subpass_description2
	pNext                   voidptr       = unsafe { nil }
	flags                   SubpassDescriptionFlags
	pipelineBindPoint       PipelineBindPoint
	viewMask                u32
	inputAttachmentCount    u32
	pInputAttachments       &AttachmentReference2
	colorAttachmentCount    u32
	pColorAttachments       &AttachmentReference2
	pResolveAttachments     &AttachmentReference2
	pDepthStencilAttachment &AttachmentReference2
	preserveAttachmentCount u32
	pPreserveAttachments    &u32
}

pub type SubpassDependency2 = C.VkSubpassDependency2

@[typedef]
pub struct C.VkSubpassDependency2 {
pub mut:
	sType           StructureType = StructureType.subpass_dependency2
	pNext           voidptr       = unsafe { nil }
	srcSubpass      u32
	dstSubpass      u32
	srcStageMask    PipelineStageFlags
	dstStageMask    PipelineStageFlags
	srcAccessMask   AccessFlags
	dstAccessMask   AccessFlags
	dependencyFlags DependencyFlags
	viewOffset      i32
}

pub type RenderPassCreateInfo2 = C.VkRenderPassCreateInfo2

@[typedef]
pub struct C.VkRenderPassCreateInfo2 {
pub mut:
	sType                   StructureType = StructureType.render_pass_create_info2
	pNext                   voidptr       = unsafe { nil }
	flags                   RenderPassCreateFlags
	attachmentCount         u32
	pAttachments            &AttachmentDescription2
	subpassCount            u32
	pSubpasses              &SubpassDescription2
	dependencyCount         u32
	pDependencies           &SubpassDependency2
	correlatedViewMaskCount u32
	pCorrelatedViewMasks    &u32
}

pub type SubpassBeginInfo = C.VkSubpassBeginInfo

@[typedef]
pub struct C.VkSubpassBeginInfo {
pub mut:
	sType    StructureType = StructureType.subpass_begin_info
	pNext    voidptr       = unsafe { nil }
	contents SubpassContents
}

pub type SubpassEndInfo = C.VkSubpassEndInfo

@[typedef]
pub struct C.VkSubpassEndInfo {
pub mut:
	sType StructureType = StructureType.subpass_end_info
	pNext voidptr       = unsafe { nil }
}

// SubpassDescriptionDepthStencilResolve extends VkSubpassDescription2
pub type SubpassDescriptionDepthStencilResolve = C.VkSubpassDescriptionDepthStencilResolve

@[typedef]
pub struct C.VkSubpassDescriptionDepthStencilResolve {
pub mut:
	sType                          StructureType = StructureType.subpass_description_depth_stencil_resolve
	pNext                          voidptr       = unsafe { nil }
	depthResolveMode               ResolveModeFlagBits
	stencilResolveMode             ResolveModeFlagBits
	pDepthStencilResolveAttachment &AttachmentReference2
}

// PhysicalDeviceDepthStencilResolveProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceDepthStencilResolveProperties = C.VkPhysicalDeviceDepthStencilResolveProperties

@[typedef]
pub struct C.VkPhysicalDeviceDepthStencilResolveProperties {
pub mut:
	sType                        StructureType = StructureType.physical_device_depth_stencil_resolve_properties
	pNext                        voidptr       = unsafe { nil }
	supportedDepthResolveModes   ResolveModeFlags
	supportedStencilResolveModes ResolveModeFlags
	independentResolveNone       Bool32
	independentResolve           Bool32
}

// ImageStencilUsageCreateInfo extends VkImageCreateInfo,VkPhysicalDeviceImageFormatInfo2
pub type ImageStencilUsageCreateInfo = C.VkImageStencilUsageCreateInfo

@[typedef]
pub struct C.VkImageStencilUsageCreateInfo {
pub mut:
	sType        StructureType = StructureType.image_stencil_usage_create_info
	pNext        voidptr       = unsafe { nil }
	stencilUsage ImageUsageFlags
}

// PhysicalDeviceImagelessFramebufferFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceImagelessFramebufferFeatures = C.VkPhysicalDeviceImagelessFramebufferFeatures

@[typedef]
pub struct C.VkPhysicalDeviceImagelessFramebufferFeatures {
pub mut:
	sType                StructureType = StructureType.physical_device_imageless_framebuffer_features
	pNext                voidptr       = unsafe { nil }
	imagelessFramebuffer Bool32
}

pub type FramebufferAttachmentImageInfo = C.VkFramebufferAttachmentImageInfo

@[typedef]
pub struct C.VkFramebufferAttachmentImageInfo {
pub mut:
	sType           StructureType = StructureType.framebuffer_attachment_image_info
	pNext           voidptr       = unsafe { nil }
	flags           ImageCreateFlags
	usage           ImageUsageFlags
	width           u32
	height          u32
	layerCount      u32
	viewFormatCount u32
	pViewFormats    &Format
}

// FramebufferAttachmentsCreateInfo extends VkFramebufferCreateInfo
pub type FramebufferAttachmentsCreateInfo = C.VkFramebufferAttachmentsCreateInfo

@[typedef]
pub struct C.VkFramebufferAttachmentsCreateInfo {
pub mut:
	sType                    StructureType = StructureType.framebuffer_attachments_create_info
	pNext                    voidptr       = unsafe { nil }
	attachmentImageInfoCount u32
	pAttachmentImageInfos    &FramebufferAttachmentImageInfo
}

// RenderPassAttachmentBeginInfo extends VkRenderPassBeginInfo
pub type RenderPassAttachmentBeginInfo = C.VkRenderPassAttachmentBeginInfo

@[typedef]
pub struct C.VkRenderPassAttachmentBeginInfo {
pub mut:
	sType           StructureType = StructureType.render_pass_attachment_begin_info
	pNext           voidptr       = unsafe { nil }
	attachmentCount u32
	pAttachments    &ImageView
}

// PhysicalDeviceSeparateDepthStencilLayoutsFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceSeparateDepthStencilLayoutsFeatures = C.VkPhysicalDeviceSeparateDepthStencilLayoutsFeatures

@[typedef]
pub struct C.VkPhysicalDeviceSeparateDepthStencilLayoutsFeatures {
pub mut:
	sType                       StructureType = StructureType.physical_device_separate_depth_stencil_layouts_features
	pNext                       voidptr       = unsafe { nil }
	separateDepthStencilLayouts Bool32
}

// AttachmentReferenceStencilLayout extends VkAttachmentReference2
pub type AttachmentReferenceStencilLayout = C.VkAttachmentReferenceStencilLayout

@[typedef]
pub struct C.VkAttachmentReferenceStencilLayout {
pub mut:
	sType         StructureType = StructureType.attachment_reference_stencil_layout
	pNext         voidptr       = unsafe { nil }
	stencilLayout ImageLayout
}

// AttachmentDescriptionStencilLayout extends VkAttachmentDescription2
pub type AttachmentDescriptionStencilLayout = C.VkAttachmentDescriptionStencilLayout

@[typedef]
pub struct C.VkAttachmentDescriptionStencilLayout {
pub mut:
	sType                StructureType = StructureType.attachment_description_stencil_layout
	pNext                voidptr       = unsafe { nil }
	stencilInitialLayout ImageLayout
	stencilFinalLayout   ImageLayout
}

@[keep_args_alive]
fn C.vkResetQueryPool(device Device, query_pool QueryPool, first_query u32, query_count u32)

pub type PFN_vkResetQueryPool = fn (device Device, query_pool QueryPool, first_query u32, query_count u32)

@[inline]
pub fn reset_query_pool(device Device,
	query_pool QueryPool,
	first_query u32,
	query_count u32) {
	C.vkResetQueryPool(device, query_pool, first_query, query_count)
}

@[keep_args_alive]
fn C.vkGetSemaphoreCounterValue(device Device, semaphore Semaphore, p_value &u64) Result

pub type PFN_vkGetSemaphoreCounterValue = fn (device Device, semaphore Semaphore, p_value &u64) Result

@[inline]
pub fn get_semaphore_counter_value(device Device,
	semaphore Semaphore,
	p_value &u64) Result {
	return C.vkGetSemaphoreCounterValue(device, semaphore, p_value)
}

@[keep_args_alive]
fn C.vkWaitSemaphores(device Device, p_wait_info &SemaphoreWaitInfo, timeout u64) Result

pub type PFN_vkWaitSemaphores = fn (device Device, p_wait_info &SemaphoreWaitInfo, timeout u64) Result

@[inline]
pub fn wait_semaphores(device Device,
	p_wait_info &SemaphoreWaitInfo,
	timeout u64) Result {
	return C.vkWaitSemaphores(device, p_wait_info, timeout)
}

@[keep_args_alive]
fn C.vkSignalSemaphore(device Device, p_signal_info &SemaphoreSignalInfo) Result

pub type PFN_vkSignalSemaphore = fn (device Device, p_signal_info &SemaphoreSignalInfo) Result

@[inline]
pub fn signal_semaphore(device Device,
	p_signal_info &SemaphoreSignalInfo) Result {
	return C.vkSignalSemaphore(device, p_signal_info)
}

@[keep_args_alive]
fn C.vkGetBufferDeviceAddress(device Device, p_info &BufferDeviceAddressInfo) DeviceAddress

pub type PFN_vkGetBufferDeviceAddress = fn (device Device, p_info &BufferDeviceAddressInfo) DeviceAddress

@[inline]
pub fn get_buffer_device_address(device Device,
	p_info &BufferDeviceAddressInfo) DeviceAddress {
	return C.vkGetBufferDeviceAddress(device, p_info)
}

@[keep_args_alive]
fn C.vkGetBufferOpaqueCaptureAddress(device Device, p_info &BufferDeviceAddressInfo) u64

pub type PFN_vkGetBufferOpaqueCaptureAddress = fn (device Device, p_info &BufferDeviceAddressInfo) u64

@[inline]
pub fn get_buffer_opaque_capture_address(device Device,
	p_info &BufferDeviceAddressInfo) u64 {
	return C.vkGetBufferOpaqueCaptureAddress(device, p_info)
}

@[keep_args_alive]
fn C.vkGetDeviceMemoryOpaqueCaptureAddress(device Device, p_info &DeviceMemoryOpaqueCaptureAddressInfo) u64

pub type PFN_vkGetDeviceMemoryOpaqueCaptureAddress = fn (device Device, p_info &DeviceMemoryOpaqueCaptureAddressInfo) u64

@[inline]
pub fn get_device_memory_opaque_capture_address(device Device,
	p_info &DeviceMemoryOpaqueCaptureAddressInfo) u64 {
	return C.vkGetDeviceMemoryOpaqueCaptureAddress(device, p_info)
}

@[keep_args_alive]
fn C.vkCmdDrawIndirectCount(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

pub type PFN_vkCmdDrawIndirectCount = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_indirect_count(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	count_buffer Buffer,
	count_buffer_offset DeviceSize,
	max_draw_count u32,
	stride u32) {
	C.vkCmdDrawIndirectCount(command_buffer, buffer, offset, count_buffer, count_buffer_offset,
		max_draw_count, stride)
}

@[keep_args_alive]
fn C.vkCmdDrawIndexedIndirectCount(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

pub type PFN_vkCmdDrawIndexedIndirectCount = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_indexed_indirect_count(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	count_buffer Buffer,
	count_buffer_offset DeviceSize,
	max_draw_count u32,
	stride u32) {
	C.vkCmdDrawIndexedIndirectCount(command_buffer, buffer, offset, count_buffer, count_buffer_offset,
		max_draw_count, stride)
}

@[keep_args_alive]
fn C.vkCreateRenderPass2(device Device, p_create_info &RenderPassCreateInfo2, p_allocator &AllocationCallbacks, p_render_pass &RenderPass) Result

pub type PFN_vkCreateRenderPass2 = fn (device Device, p_create_info &RenderPassCreateInfo2, p_allocator &AllocationCallbacks, p_render_pass &RenderPass) Result

@[inline]
pub fn create_render_pass2(device Device,
	p_create_info &RenderPassCreateInfo2,
	p_allocator &AllocationCallbacks,
	p_render_pass &RenderPass) Result {
	return C.vkCreateRenderPass2(device, p_create_info, p_allocator, p_render_pass)
}

@[keep_args_alive]
fn C.vkCmdBeginRenderPass2(command_buffer CommandBuffer, p_render_pass_begin &RenderPassBeginInfo, p_subpass_begin_info &SubpassBeginInfo)

pub type PFN_vkCmdBeginRenderPass2 = fn (command_buffer CommandBuffer, p_render_pass_begin &RenderPassBeginInfo, p_subpass_begin_info &SubpassBeginInfo)

@[inline]
pub fn cmd_begin_render_pass2(command_buffer CommandBuffer,
	p_render_pass_begin &RenderPassBeginInfo,
	p_subpass_begin_info &SubpassBeginInfo) {
	C.vkCmdBeginRenderPass2(command_buffer, p_render_pass_begin, p_subpass_begin_info)
}

@[keep_args_alive]
fn C.vkCmdNextSubpass2(command_buffer CommandBuffer, p_subpass_begin_info &SubpassBeginInfo, p_subpass_end_info &SubpassEndInfo)

pub type PFN_vkCmdNextSubpass2 = fn (command_buffer CommandBuffer, p_subpass_begin_info &SubpassBeginInfo, p_subpass_end_info &SubpassEndInfo)

@[inline]
pub fn cmd_next_subpass2(command_buffer CommandBuffer,
	p_subpass_begin_info &SubpassBeginInfo,
	p_subpass_end_info &SubpassEndInfo) {
	C.vkCmdNextSubpass2(command_buffer, p_subpass_begin_info, p_subpass_end_info)
}

@[keep_args_alive]
fn C.vkCmdEndRenderPass2(command_buffer CommandBuffer, p_subpass_end_info &SubpassEndInfo)

pub type PFN_vkCmdEndRenderPass2 = fn (command_buffer CommandBuffer, p_subpass_end_info &SubpassEndInfo)

@[inline]
pub fn cmd_end_render_pass2(command_buffer CommandBuffer,
	p_subpass_end_info &SubpassEndInfo) {
	C.vkCmdEndRenderPass2(command_buffer, p_subpass_end_info)
}

pub const api_version_1_3 = make_api_version(0, 1, 3, 0) // patch version should always be set to 0

pub type Flags64 = u64

// Pointer to VkPrivateDataSlot_T
pub type PrivateDataSlot = voidptr

pub enum ToolPurposeFlagBits as u32 {
	validation              = u32(0x00000001)
	profiling               = u32(0x00000002)
	tracing                 = u32(0x00000004)
	additional_features     = u32(0x00000008)
	modifying_features      = u32(0x00000010)
	debug_reporting_bit_ext = u32(0x00000020)
	debug_markers_bit_ext   = u32(0x00000040)
	max_enum                = max_int
}
pub type ToolPurposeFlags = u32
pub type PrivateDataSlotCreateFlags = u32
pub type PipelineStageFlags2 = u64

// Flag bits for PipelineStageFlagBits2
pub type PipelineStageFlagBits2 = u64

pub const pipeline_stage_2_none = u64(0)
pub const pipeline_stage_2_top_of_pipe_bit = u64(0x00000001)
pub const pipeline_stage_2_draw_indirect_bit = u64(0x00000002)
pub const pipeline_stage_2_vertex_input_bit = u64(0x00000004)
pub const pipeline_stage_2_vertex_shader_bit = u64(0x00000008)
pub const pipeline_stage_2_tessellation_control_shader_bit = u64(0x00000010)
pub const pipeline_stage_2_tessellation_evaluation_shader_bit = u64(0x00000020)
pub const pipeline_stage_2_geometry_shader_bit = u64(0x00000040)
pub const pipeline_stage_2_fragment_shader_bit = u64(0x00000080)
pub const pipeline_stage_2_early_fragment_tests_bit = u64(0x00000100)
pub const pipeline_stage_2_late_fragment_tests_bit = u64(0x00000200)
pub const pipeline_stage_2_color_attachment_output_bit = u64(0x00000400)
pub const pipeline_stage_2_compute_shader_bit = u64(0x00000800)
pub const pipeline_stage_2_all_transfer_bit = u64(0x00001000)
pub const pipeline_stage_2_transfer_bit = pipeline_stage_2_all_transfer_bit
pub const pipeline_stage_2_bottom_of_pipe_bit = u64(0x00002000)
pub const pipeline_stage_2_host_bit = u64(0x00004000)
pub const pipeline_stage_2_all_graphics_bit = u64(0x00008000)
pub const pipeline_stage_2_all_commands_bit = u64(0x00010000)
pub const pipeline_stage_2_copy_bit = u64(0x100000000)
pub const pipeline_stage_2_resolve_bit = u64(0x200000000)
pub const pipeline_stage_2_blit_bit = u64(0x400000000)
pub const pipeline_stage_2_clear_bit = u64(0x800000000)
pub const pipeline_stage_2_index_input_bit = u64(0x1000000000)
pub const pipeline_stage_2_vertex_attribute_input_bit = u64(0x2000000000)
pub const pipeline_stage_2_pre_rasterization_shaders_bit = u64(0x4000000000)
pub const pipeline_stage_2_video_decode_bit_khr = u64(0x04000000)
pub const pipeline_stage_2_video_encode_bit_khr = u64(0x08000000)
pub const pipeline_stage_2_none_khr = pipeline_stage_2_none
pub const pipeline_stage_2_top_of_pipe_bit_khr = pipeline_stage_2_top_of_pipe_bit
pub const pipeline_stage_2_draw_indirect_bit_khr = pipeline_stage_2_draw_indirect_bit
pub const pipeline_stage_2_vertex_input_bit_khr = u32(pipeline_stage_2_vertex_input_bit)
pub const pipeline_stage_2_vertex_shader_bit_khr = pipeline_stage_2_vertex_shader_bit
pub const pipeline_stage_2_tessellation_control_shader_bit_khr = pipeline_stage_2_tessellation_control_shader_bit
pub const pipeline_stage_2_tessellation_evaluation_shader_bit_khr = u32(pipeline_stage_2_tessellation_evaluation_shader_bit)
pub const pipeline_stage_2_geometry_shader_bit_khr = pipeline_stage_2_geometry_shader_bit
pub const pipeline_stage_2_fragment_shader_bit_khr = pipeline_stage_2_fragment_shader_bit
pub const pipeline_stage_2_early_fragment_tests_bit_khr = pipeline_stage_2_early_fragment_tests_bit
pub const pipeline_stage_2_late_fragment_tests_bit_khr = pipeline_stage_2_late_fragment_tests_bit
pub const pipeline_stage_2_color_attachment_output_bit_khr = u32(pipeline_stage_2_color_attachment_output_bit)
pub const pipeline_stage_2_compute_shader_bit_khr = u32(pipeline_stage_2_compute_shader_bit)
pub const pipeline_stage_2_all_transfer_bit_khr = pipeline_stage_2_all_transfer_bit
pub const pipeline_stage_2_transfer_bit_khr = pipeline_stage_2_all_transfer_bit
pub const pipeline_stage_2_bottom_of_pipe_bit_khr = pipeline_stage_2_bottom_of_pipe_bit
pub const pipeline_stage_2_host_bit_khr = pipeline_stage_2_host_bit
pub const pipeline_stage_2_all_graphics_bit_khr = pipeline_stage_2_all_graphics_bit
pub const pipeline_stage_2_all_commands_bit_khr = pipeline_stage_2_all_commands_bit
pub const pipeline_stage_2_copy_bit_khr = pipeline_stage_2_copy_bit
pub const pipeline_stage_2_resolve_bit_khr = pipeline_stage_2_resolve_bit
pub const pipeline_stage_2_blit_bit_khr = pipeline_stage_2_blit_bit
pub const pipeline_stage_2_clear_bit_khr = pipeline_stage_2_clear_bit
pub const pipeline_stage_2_index_input_bit_khr = u32(pipeline_stage_2_index_input_bit)
pub const pipeline_stage_2_vertex_attribute_input_bit_khr = u32(pipeline_stage_2_vertex_attribute_input_bit)
pub const pipeline_stage_2_pre_rasterization_shaders_bit_khr = pipeline_stage_2_pre_rasterization_shaders_bit
pub const pipeline_stage_2_transform_feedback_bit_ext = u64(0x01000000)
pub const pipeline_stage_2_conditional_rendering_bit_ext = u64(0x00040000)
pub const pipeline_stage_2_command_preprocess_bit_nv = pipeline_stage_2_command_preprocess_bit_ext
pub const pipeline_stage_2_command_preprocess_bit_ext = u64(0x00020000)
pub const pipeline_stage_2_fragment_shading_rate_attachment_bit_khr = u64(0x00400000)
pub const pipeline_stage_2_shading_rate_image_bit_nv = pipeline_stage_2_fragment_shading_rate_attachment_bit_khr
pub const pipeline_stage_2_acceleration_structure_build_bit_khr = u64(0x02000000)
pub const pipeline_stage_2_ray_tracing_shader_bit_khr = u64(0x00200000)
pub const pipeline_stage_2_ray_tracing_shader_bit_nv = pipeline_stage_2_ray_tracing_shader_bit_khr
pub const pipeline_stage_2_acceleration_structure_build_bit_nv = u32(pipeline_stage_2_acceleration_structure_build_bit_khr)
pub const pipeline_stage_2_fragment_density_process_bit_ext = u64(0x00800000)
pub const pipeline_stage_2_task_shader_bit_nv = pipeline_stage_2_task_shader_bit_ext
pub const pipeline_stage_2_mesh_shader_bit_nv = pipeline_stage_2_mesh_shader_bit_ext
pub const pipeline_stage_2_task_shader_bit_ext = u64(0x00080000)
pub const pipeline_stage_2_mesh_shader_bit_ext = u64(0x00100000)
pub const pipeline_stage_2_subpass_shader_bit_huawei = u64(0x8000000000)
// VK_PIPELINE_STAGE_2_SUBPASS_SHADING_BIT_HUAWEI is a deprecated alias
pub const pipeline_stage_2_subpass_shading_bit_huawei = u32(pipeline_stage_2_subpass_shader_bit_huawei)
pub const pipeline_stage_2_invocation_mask_bit_huawei = u64(0x10000000000)
pub const pipeline_stage_2_acceleration_structure_copy_bit_khr = u64(0x10000000)
pub const pipeline_stage_2_micromap_build_bit_ext = u64(0x40000000)
pub const pipeline_stage_2_cluster_culling_shader_bit_huawei = u64(0x20000000000)
pub const pipeline_stage_2_optical_flow_bit_nv = u64(0x20000000)
pub const pipeline_stage_2_convert_cooperative_vector_matrix_bit_nv = u64(0x100000000000)
pub const pipeline_stage_2_data_graph_bit_arm = u64(0x40000000000)
pub const pipeline_stage_2_copy_indirect_bit_khr = u64(0x400000000000)
pub const pipeline_stage_2_memory_decompression_bit_ext = u64(0x200000000000)

pub type AccessFlags2 = u64

// Flag bits for AccessFlagBits2
pub type AccessFlagBits2 = u64

pub const access_2_none = u64(0)
pub const access_2_indirect_command_read_bit = u64(0x00000001)
pub const access_2_index_read_bit = u64(0x00000002)
pub const access_2_vertex_attribute_read_bit = u64(0x00000004)
pub const access_2_uniform_read_bit = u64(0x00000008)
pub const access_2_input_attachment_read_bit = u64(0x00000010)
pub const access_2_shader_read_bit = u64(0x00000020)
pub const access_2_shader_write_bit = u64(0x00000040)
pub const access_2_color_attachment_read_bit = u64(0x00000080)
pub const access_2_color_attachment_write_bit = u64(0x00000100)
pub const access_2_depth_stencil_attachment_read_bit = u64(0x00000200)
pub const access_2_depth_stencil_attachment_write_bit = u64(0x00000400)
pub const access_2_transfer_read_bit = u64(0x00000800)
pub const access_2_transfer_write_bit = u64(0x00001000)
pub const access_2_host_read_bit = u64(0x00002000)
pub const access_2_host_write_bit = u64(0x00004000)
pub const access_2_memory_read_bit = u64(0x00008000)
pub const access_2_memory_write_bit = u64(0x00010000)
pub const access_2_shader_sampled_read_bit = u64(0x100000000)
pub const access_2_shader_storage_read_bit = u64(0x200000000)
pub const access_2_shader_storage_write_bit = u64(0x400000000)
pub const access_2_video_decode_read_bit_khr = u64(0x800000000)
pub const access_2_video_decode_write_bit_khr = u64(0x1000000000)
pub const access_2_video_encode_read_bit_khr = u64(0x2000000000)
pub const access_2_video_encode_write_bit_khr = u64(0x4000000000)
pub const access_2_shader_tile_attachment_read_bit_qcom = u64(0x8000000000000)
pub const access_2_shader_tile_attachment_write_bit_qcom = u64(0x10000000000000)
pub const access_2_none_khr = access_2_none
pub const access_2_indirect_command_read_bit_khr = access_2_indirect_command_read_bit
pub const access_2_index_read_bit_khr = access_2_index_read_bit
pub const access_2_vertex_attribute_read_bit_khr = u32(access_2_vertex_attribute_read_bit)
pub const access_2_uniform_read_bit_khr = u32(access_2_uniform_read_bit)
pub const access_2_input_attachment_read_bit_khr = u32(access_2_input_attachment_read_bit)
pub const access_2_shader_read_bit_khr = access_2_shader_read_bit
pub const access_2_shader_write_bit_khr = access_2_shader_write_bit
pub const access_2_color_attachment_read_bit_khr = access_2_color_attachment_read_bit
pub const access_2_color_attachment_write_bit_khr = access_2_color_attachment_write_bit
pub const access_2_depth_stencil_attachment_read_bit_khr = access_2_depth_stencil_attachment_read_bit
pub const access_2_depth_stencil_attachment_write_bit_khr = access_2_depth_stencil_attachment_write_bit
pub const access_2_transfer_read_bit_khr = access_2_transfer_read_bit
pub const access_2_transfer_write_bit_khr = access_2_transfer_write_bit
pub const access_2_host_read_bit_khr = access_2_host_read_bit
pub const access_2_host_write_bit_khr = access_2_host_write_bit
pub const access_2_memory_read_bit_khr = access_2_memory_read_bit
pub const access_2_memory_write_bit_khr = access_2_memory_write_bit
pub const access_2_shader_sampled_read_bit_khr = access_2_shader_sampled_read_bit
pub const access_2_shader_storage_read_bit_khr = access_2_shader_storage_read_bit
pub const access_2_shader_storage_write_bit_khr = access_2_shader_storage_write_bit
pub const access_2_transform_feedback_write_bit_ext = u64(0x02000000)
pub const access_2_transform_feedback_counter_read_bit_ext = u64(0x04000000)
pub const access_2_transform_feedback_counter_write_bit_ext = u64(0x08000000)
pub const access_2_conditional_rendering_read_bit_ext = u64(0x00100000)
pub const access_2_command_preprocess_read_bit_nv = access_2_command_preprocess_read_bit_ext
pub const access_2_command_preprocess_write_bit_nv = access_2_command_preprocess_write_bit_ext
pub const access_2_command_preprocess_read_bit_ext = u64(0x00020000)
pub const access_2_command_preprocess_write_bit_ext = u64(0x00040000)
pub const access_2_fragment_shading_rate_attachment_read_bit_khr = u64(0x00800000)
pub const access_2_shading_rate_image_read_bit_nv = access_2_fragment_shading_rate_attachment_read_bit_khr
pub const access_2_acceleration_structure_read_bit_khr = u64(0x00200000)
pub const access_2_acceleration_structure_write_bit_khr = u64(0x00400000)
pub const access_2_acceleration_structure_read_bit_nv = u32(access_2_acceleration_structure_read_bit_khr)
pub const access_2_acceleration_structure_write_bit_nv = u32(access_2_acceleration_structure_write_bit_khr)
pub const access_2_fragment_density_map_read_bit_ext = u64(0x01000000)
pub const access_2_color_attachment_read_noncoherent_bit_ext = u64(0x00080000)
pub const access_2_descriptor_buffer_read_bit_ext = u64(0x20000000000)
pub const access_2_invocation_mask_read_bit_huawei = u64(0x8000000000)
pub const access_2_shader_binding_table_read_bit_khr = u64(0x10000000000)
pub const access_2_micromap_read_bit_ext = u64(0x100000000000)
pub const access_2_micromap_write_bit_ext = u64(0x200000000000)
pub const access_2_optical_flow_read_bit_nv = u64(0x40000000000)
pub const access_2_optical_flow_write_bit_nv = u64(0x80000000000)
pub const access_2_data_graph_read_bit_arm = u64(0x800000000000)
pub const access_2_data_graph_write_bit_arm = u64(0x1000000000000)
pub const access_2_memory_decompression_read_bit_ext = u64(0x80000000000000)
pub const access_2_memory_decompression_write_bit_ext = u64(0x100000000000000)

pub enum SubmitFlagBits as u32 {
	protected = u32(0x00000001)
	max_enum  = max_int
}
pub type SubmitFlags = u32
pub type FormatFeatureFlags2 = u64

// Flag bits for FormatFeatureFlagBits2
pub type FormatFeatureFlagBits2 = u64

pub const format_feature_2_sampled_image_bit = u64(0x00000001)
pub const format_feature_2_storage_image_bit = u64(0x00000002)
pub const format_feature_2_storage_image_atomic_bit = u64(0x00000004)
pub const format_feature_2_uniform_texel_buffer_bit = u64(0x00000008)
pub const format_feature_2_storage_texel_buffer_bit = u64(0x00000010)
pub const format_feature_2_storage_texel_buffer_atomic_bit = u64(0x00000020)
pub const format_feature_2_vertex_buffer_bit = u64(0x00000040)
pub const format_feature_2_color_attachment_bit = u64(0x00000080)
pub const format_feature_2_color_attachment_blend_bit = u64(0x00000100)
pub const format_feature_2_depth_stencil_attachment_bit = u64(0x00000200)
pub const format_feature_2_blit_src_bit = u64(0x00000400)
pub const format_feature_2_blit_dst_bit = u64(0x00000800)
pub const format_feature_2_sampled_image_filter_linear_bit = u64(0x00001000)
pub const format_feature_2_transfer_src_bit = u64(0x00004000)
pub const format_feature_2_transfer_dst_bit = u64(0x00008000)
pub const format_feature_2_sampled_image_filter_minmax_bit = u64(0x00010000)
pub const format_feature_2_midpoint_chroma_samples_bit = u64(0x00020000)
pub const format_feature_2_sampled_image_ycbcr_conversion_linear_filter_bit = u64(0x00040000)
pub const format_feature_2_sampled_image_ycbcr_conversion_separate_reconstruction_filter_bit = u64(0x00080000)
pub const format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_bit = u64(0x00100000)
pub const format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_forceable_bit = u64(0x00200000)
pub const format_feature_2_disjoint_bit = u64(0x00400000)
pub const format_feature_2_cosited_chroma_samples_bit = u64(0x00800000)
pub const format_feature_2_storage_read_without_format_bit = u64(0x80000000)
pub const format_feature_2_storage_write_without_format_bit = u64(0x100000000)
pub const format_feature_2_sampled_image_depth_comparison_bit = u64(0x200000000)
pub const format_feature_2_sampled_image_filter_cubic_bit = u64(0x00002000)
pub const format_feature_2_host_image_transfer_bit = u64(0x400000000000)
pub const format_feature_2_video_decode_output_bit_khr = u64(0x02000000)
pub const format_feature_2_video_decode_dpb_bit_khr = u64(0x04000000)
pub const format_feature_2_acceleration_structure_vertex_buffer_bit_khr = u64(0x20000000)
pub const format_feature_2_fragment_density_map_bit_ext = u64(0x01000000)
pub const format_feature_2_fragment_shading_rate_attachment_bit_khr = u64(0x40000000)
pub const format_feature_2_host_image_transfer_bit_ext = u32(format_feature_2_host_image_transfer_bit)
pub const format_feature_2_video_encode_input_bit_khr = u64(0x08000000)
pub const format_feature_2_video_encode_dpb_bit_khr = u64(0x10000000)
pub const format_feature_2_sampled_image_bit_khr = u32(format_feature_2_sampled_image_bit)
pub const format_feature_2_storage_image_bit_khr = u32(format_feature_2_storage_image_bit)
pub const format_feature_2_storage_image_atomic_bit_khr = u32(format_feature_2_storage_image_atomic_bit)
pub const format_feature_2_uniform_texel_buffer_bit_khr = u32(format_feature_2_uniform_texel_buffer_bit)
pub const format_feature_2_storage_texel_buffer_bit_khr = u32(format_feature_2_storage_texel_buffer_bit)
pub const format_feature_2_storage_texel_buffer_atomic_bit_khr = u32(format_feature_2_storage_texel_buffer_atomic_bit)
pub const format_feature_2_vertex_buffer_bit_khr = u32(format_feature_2_vertex_buffer_bit)
pub const format_feature_2_color_attachment_bit_khr = u32(format_feature_2_color_attachment_bit)
pub const format_feature_2_color_attachment_blend_bit_khr = u32(format_feature_2_color_attachment_blend_bit)
pub const format_feature_2_depth_stencil_attachment_bit_khr = u32(format_feature_2_depth_stencil_attachment_bit)
pub const format_feature_2_blit_src_bit_khr = u32(format_feature_2_blit_src_bit)
pub const format_feature_2_blit_dst_bit_khr = u32(format_feature_2_blit_dst_bit)
pub const format_feature_2_sampled_image_filter_linear_bit_khr = u32(format_feature_2_sampled_image_filter_linear_bit)
pub const format_feature_2_transfer_src_bit_khr = u32(format_feature_2_transfer_src_bit)
pub const format_feature_2_transfer_dst_bit_khr = u32(format_feature_2_transfer_dst_bit)
pub const format_feature_2_midpoint_chroma_samples_bit_khr = u32(format_feature_2_midpoint_chroma_samples_bit)
pub const format_feature_2_sampled_image_ycbcr_conversion_linear_filter_bit_khr = u32(format_feature_2_sampled_image_ycbcr_conversion_linear_filter_bit)
pub const format_feature_2_sampled_image_ycbcr_conversion_separate_reconstruction_filter_bit_khr = u32(format_feature_2_sampled_image_ycbcr_conversion_separate_reconstruction_filter_bit)
pub const format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_bit_khr = u32(format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_bit)
pub const format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_forceable_bit_khr = u32(format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_forceable_bit)
pub const format_feature_2_disjoint_bit_khr = u32(format_feature_2_disjoint_bit)
pub const format_feature_2_cosited_chroma_samples_bit_khr = u32(format_feature_2_cosited_chroma_samples_bit)
pub const format_feature_2_storage_read_without_format_bit_khr = u32(format_feature_2_storage_read_without_format_bit)
pub const format_feature_2_storage_write_without_format_bit_khr = u32(format_feature_2_storage_write_without_format_bit)
pub const format_feature_2_sampled_image_depth_comparison_bit_khr = u32(format_feature_2_sampled_image_depth_comparison_bit)
pub const format_feature_2_sampled_image_filter_minmax_bit_khr = u32(format_feature_2_sampled_image_filter_minmax_bit)
pub const format_feature_2_sampled_image_filter_cubic_bit_ext = u32(format_feature_2_sampled_image_filter_cubic_bit)
pub const format_feature_2_acceleration_structure_radius_buffer_bit_nv = u64(0x8000000000000)
pub const format_feature_2_linear_color_attachment_bit_nv = u64(0x4000000000)
pub const format_feature_2_weight_image_bit_qcom = u64(0x400000000)
pub const format_feature_2_weight_sampled_image_bit_qcom = u64(0x800000000)
pub const format_feature_2_block_matching_bit_qcom = u64(0x1000000000)
pub const format_feature_2_box_filter_sampled_bit_qcom = u64(0x2000000000)
pub const format_feature_2_tensor_shader_bit_arm = u64(0x8000000000)
pub const format_feature_2_tensor_image_aliasing_bit_arm = u64(0x80000000000)
pub const format_feature_2_optical_flow_image_bit_nv = u64(0x10000000000)
pub const format_feature_2_optical_flow_vector_bit_nv = u64(0x20000000000)
pub const format_feature_2_optical_flow_cost_bit_nv = u64(0x40000000000)
pub const format_feature_2_tensor_data_graph_bit_arm = u64(0x1000000000000)
pub const format_feature_2_copy_image_indirect_dst_bit_khr = u64(0x800000000000000)
pub const format_feature_2_video_encode_quantization_delta_map_bit_khr = u64(0x2000000000000)
pub const format_feature_2_video_encode_emphasis_map_bit_khr = u64(0x4000000000000)
pub const format_feature_2_depth_copy_on_compute_queue_bit_khr = u64(0x10000000000000)
pub const format_feature_2_depth_copy_on_transfer_queue_bit_khr = u64(0x20000000000000)
pub const format_feature_2_stencil_copy_on_compute_queue_bit_khr = u64(0x40000000000000)
pub const format_feature_2_stencil_copy_on_transfer_queue_bit_khr = u64(0x80000000000000)

pub enum PipelineCreationFeedbackFlagBits as u32 {
	valid                          = u32(0x00000001)
	application_pipeline_cache_hit = u32(0x00000002)
	base_pipeline_acceleration     = u32(0x00000004)
	max_enum                       = max_int
}
pub type PipelineCreationFeedbackFlags = u32

pub enum RenderingFlagBits as u32 {
	contents_secondary_command_buffers   = u32(0x00000001)
	suspending                           = u32(0x00000002)
	resuming                             = u32(0x00000004)
	enable_legacy_dithering_bit_ext      = u32(0x00000008)
	contents_inline                      = u32(0x00000010)
	per_layer_fragment_density_bit_valve = u32(0x00000020)
	local_read_concurrent_access_control = u32(0x00000100)
	max_enum                             = max_int
}
pub type RenderingFlags = u32

// PhysicalDeviceVulkan13Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVulkan13Features = C.VkPhysicalDeviceVulkan13Features

@[typedef]
pub struct C.VkPhysicalDeviceVulkan13Features {
pub mut:
	sType                                              StructureType = StructureType.physical_device_vulkan1_3_features
	pNext                                              voidptr       = unsafe { nil }
	robustImageAccess                                  Bool32
	inlineUniformBlock                                 Bool32
	descriptorBindingInlineUniformBlockUpdateAfterBind Bool32
	pipelineCreationCacheControl                       Bool32
	privateData                                        Bool32
	shaderDemoteToHelperInvocation                     Bool32
	shaderTerminateInvocation                          Bool32
	subgroupSizeControl                                Bool32
	computeFullSubgroups                               Bool32
	synchronization2                                   Bool32
	textureCompressionASTC_HDR                         Bool32
	shaderZeroInitializeWorkgroupMemory                Bool32
	dynamicRendering                                   Bool32
	shaderIntegerDotProduct                            Bool32
	maintenance4                                       Bool32
}

// PhysicalDeviceVulkan13Properties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceVulkan13Properties = C.VkPhysicalDeviceVulkan13Properties

@[typedef]
pub struct C.VkPhysicalDeviceVulkan13Properties {
pub mut:
	sType                                                                         StructureType = StructureType.physical_device_vulkan1_3_properties
	pNext                                                                         voidptr       = unsafe { nil }
	minSubgroupSize                                                               u32
	maxSubgroupSize                                                               u32
	maxComputeWorkgroupSubgroups                                                  u32
	requiredSubgroupSizeStages                                                    ShaderStageFlags
	maxInlineUniformBlockSize                                                     u32
	maxPerStageDescriptorInlineUniformBlocks                                      u32
	maxPerStageDescriptorUpdateAfterBindInlineUniformBlocks                       u32
	maxDescriptorSetInlineUniformBlocks                                           u32
	maxDescriptorSetUpdateAfterBindInlineUniformBlocks                            u32
	maxInlineUniformTotalSize                                                     u32
	integerDotProduct8BitUnsignedAccelerated                                      Bool32
	integerDotProduct8BitSignedAccelerated                                        Bool32
	integerDotProduct8BitMixedSignednessAccelerated                               Bool32
	integerDotProduct4x8BitPackedUnsignedAccelerated                              Bool32
	integerDotProduct4x8BitPackedSignedAccelerated                                Bool32
	integerDotProduct4x8BitPackedMixedSignednessAccelerated                       Bool32
	integerDotProduct16BitUnsignedAccelerated                                     Bool32
	integerDotProduct16BitSignedAccelerated                                       Bool32
	integerDotProduct16BitMixedSignednessAccelerated                              Bool32
	integerDotProduct32BitUnsignedAccelerated                                     Bool32
	integerDotProduct32BitSignedAccelerated                                       Bool32
	integerDotProduct32BitMixedSignednessAccelerated                              Bool32
	integerDotProduct64BitUnsignedAccelerated                                     Bool32
	integerDotProduct64BitSignedAccelerated                                       Bool32
	integerDotProduct64BitMixedSignednessAccelerated                              Bool32
	integerDotProductAccumulatingSaturating8BitUnsignedAccelerated                Bool32
	integerDotProductAccumulatingSaturating8BitSignedAccelerated                  Bool32
	integerDotProductAccumulatingSaturating8BitMixedSignednessAccelerated         Bool32
	integerDotProductAccumulatingSaturating4x8BitPackedUnsignedAccelerated        Bool32
	integerDotProductAccumulatingSaturating4x8BitPackedSignedAccelerated          Bool32
	integerDotProductAccumulatingSaturating4x8BitPackedMixedSignednessAccelerated Bool32
	integerDotProductAccumulatingSaturating16BitUnsignedAccelerated               Bool32
	integerDotProductAccumulatingSaturating16BitSignedAccelerated                 Bool32
	integerDotProductAccumulatingSaturating16BitMixedSignednessAccelerated        Bool32
	integerDotProductAccumulatingSaturating32BitUnsignedAccelerated               Bool32
	integerDotProductAccumulatingSaturating32BitSignedAccelerated                 Bool32
	integerDotProductAccumulatingSaturating32BitMixedSignednessAccelerated        Bool32
	integerDotProductAccumulatingSaturating64BitUnsignedAccelerated               Bool32
	integerDotProductAccumulatingSaturating64BitSignedAccelerated                 Bool32
	integerDotProductAccumulatingSaturating64BitMixedSignednessAccelerated        Bool32
	storageTexelBufferOffsetAlignmentBytes                                        DeviceSize
	storageTexelBufferOffsetSingleTexelAlignment                                  Bool32
	uniformTexelBufferOffsetAlignmentBytes                                        DeviceSize
	uniformTexelBufferOffsetSingleTexelAlignment                                  Bool32
	maxBufferSize                                                                 DeviceSize
}

pub type PhysicalDeviceToolProperties = C.VkPhysicalDeviceToolProperties

@[typedef]
pub struct C.VkPhysicalDeviceToolProperties {
pub mut:
	sType       StructureType = StructureType.physical_device_tool_properties
	pNext       voidptr       = unsafe { nil }
	name        [max_extension_name_size]char
	version     [max_extension_name_size]char
	purposes    ToolPurposeFlags
	description [max_description_size]char
	layer       [max_extension_name_size]char
}

// PhysicalDevicePrivateDataFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePrivateDataFeatures = C.VkPhysicalDevicePrivateDataFeatures

@[typedef]
pub struct C.VkPhysicalDevicePrivateDataFeatures {
pub mut:
	sType       StructureType = StructureType.physical_device_private_data_features
	pNext       voidptr       = unsafe { nil }
	privateData Bool32
}

// DevicePrivateDataCreateInfo extends VkDeviceCreateInfo
pub type DevicePrivateDataCreateInfo = C.VkDevicePrivateDataCreateInfo

@[typedef]
pub struct C.VkDevicePrivateDataCreateInfo {
pub mut:
	sType                       StructureType = StructureType.device_private_data_create_info
	pNext                       voidptr       = unsafe { nil }
	privateDataSlotRequestCount u32
}

pub type PrivateDataSlotCreateInfo = C.VkPrivateDataSlotCreateInfo

@[typedef]
pub struct C.VkPrivateDataSlotCreateInfo {
pub mut:
	sType StructureType = StructureType.private_data_slot_create_info
	pNext voidptr       = unsafe { nil }
	flags PrivateDataSlotCreateFlags
}

// MemoryBarrier2 extends VkSubpassDependency2
pub type MemoryBarrier2 = C.VkMemoryBarrier2

@[typedef]
pub struct C.VkMemoryBarrier2 {
pub mut:
	sType         StructureType = StructureType.memory_barrier2
	pNext         voidptr       = unsafe { nil }
	srcStageMask  PipelineStageFlags2
	srcAccessMask AccessFlags2
	dstStageMask  PipelineStageFlags2
	dstAccessMask AccessFlags2
}

pub type BufferMemoryBarrier2 = C.VkBufferMemoryBarrier2

@[typedef]
pub struct C.VkBufferMemoryBarrier2 {
pub mut:
	sType               StructureType = StructureType.buffer_memory_barrier2
	pNext               voidptr       = unsafe { nil }
	srcStageMask        PipelineStageFlags2
	srcAccessMask       AccessFlags2
	dstStageMask        PipelineStageFlags2
	dstAccessMask       AccessFlags2
	srcQueueFamilyIndex u32
	dstQueueFamilyIndex u32
	buffer              Buffer
	offset              DeviceSize
	size                DeviceSize
}

pub type ImageMemoryBarrier2 = C.VkImageMemoryBarrier2

@[typedef]
pub struct C.VkImageMemoryBarrier2 {
pub mut:
	sType               StructureType = StructureType.image_memory_barrier2
	pNext               voidptr       = unsafe { nil }
	srcStageMask        PipelineStageFlags2
	srcAccessMask       AccessFlags2
	dstStageMask        PipelineStageFlags2
	dstAccessMask       AccessFlags2
	oldLayout           ImageLayout
	newLayout           ImageLayout
	srcQueueFamilyIndex u32
	dstQueueFamilyIndex u32
	image               Image
	subresourceRange    ImageSubresourceRange
}

pub type DependencyInfo = C.VkDependencyInfo

@[typedef]
pub struct C.VkDependencyInfo {
pub mut:
	sType                    StructureType = StructureType.dependency_info
	pNext                    voidptr       = unsafe { nil }
	dependencyFlags          DependencyFlags
	memoryBarrierCount       u32
	pMemoryBarriers          &MemoryBarrier2
	bufferMemoryBarrierCount u32
	pBufferMemoryBarriers    &BufferMemoryBarrier2
	imageMemoryBarrierCount  u32
	pImageMemoryBarriers     &ImageMemoryBarrier2
}

pub type SemaphoreSubmitInfo = C.VkSemaphoreSubmitInfo

@[typedef]
pub struct C.VkSemaphoreSubmitInfo {
pub mut:
	sType       StructureType = StructureType.semaphore_submit_info
	pNext       voidptr       = unsafe { nil }
	semaphore   Semaphore
	value       u64
	stageMask   PipelineStageFlags2
	deviceIndex u32
}

pub type CommandBufferSubmitInfo = C.VkCommandBufferSubmitInfo

@[typedef]
pub struct C.VkCommandBufferSubmitInfo {
pub mut:
	sType         StructureType = StructureType.command_buffer_submit_info
	pNext         voidptr       = unsafe { nil }
	commandBuffer CommandBuffer
	deviceMask    u32
}

pub type SubmitInfo2 = C.VkSubmitInfo2

@[typedef]
pub struct C.VkSubmitInfo2 {
pub mut:
	sType                    StructureType = StructureType.submit_info2
	pNext                    voidptr       = unsafe { nil }
	flags                    SubmitFlags
	waitSemaphoreInfoCount   u32
	pWaitSemaphoreInfos      &SemaphoreSubmitInfo
	commandBufferInfoCount   u32
	pCommandBufferInfos      &CommandBufferSubmitInfo
	signalSemaphoreInfoCount u32
	pSignalSemaphoreInfos    &SemaphoreSubmitInfo
}

// PhysicalDeviceSynchronization2Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceSynchronization2Features = C.VkPhysicalDeviceSynchronization2Features

@[typedef]
pub struct C.VkPhysicalDeviceSynchronization2Features {
pub mut:
	sType            StructureType = StructureType.physical_device_synchronization2_features
	pNext            voidptr       = unsafe { nil }
	synchronization2 Bool32
}

pub type BufferCopy2 = C.VkBufferCopy2

@[typedef]
pub struct C.VkBufferCopy2 {
pub mut:
	sType     StructureType = StructureType.buffer_copy2
	pNext     voidptr       = unsafe { nil }
	srcOffset DeviceSize
	dstOffset DeviceSize
	size      DeviceSize
}

pub type CopyBufferInfo2 = C.VkCopyBufferInfo2

@[typedef]
pub struct C.VkCopyBufferInfo2 {
pub mut:
	sType       StructureType = StructureType.copy_buffer_info2
	pNext       voidptr       = unsafe { nil }
	srcBuffer   Buffer
	dstBuffer   Buffer
	regionCount u32
	pRegions    &BufferCopy2
}

pub type ImageCopy2 = C.VkImageCopy2

@[typedef]
pub struct C.VkImageCopy2 {
pub mut:
	sType          StructureType = StructureType.image_copy2
	pNext          voidptr       = unsafe { nil }
	srcSubresource ImageSubresourceLayers
	srcOffset      Offset3D
	dstSubresource ImageSubresourceLayers
	dstOffset      Offset3D
	extent         Extent3D
}

pub type CopyImageInfo2 = C.VkCopyImageInfo2

@[typedef]
pub struct C.VkCopyImageInfo2 {
pub mut:
	sType          StructureType = StructureType.copy_image_info2
	pNext          voidptr       = unsafe { nil }
	srcImage       Image
	srcImageLayout ImageLayout
	dstImage       Image
	dstImageLayout ImageLayout
	regionCount    u32
	pRegions       &ImageCopy2
}

pub type BufferImageCopy2 = C.VkBufferImageCopy2

@[typedef]
pub struct C.VkBufferImageCopy2 {
pub mut:
	sType             StructureType = StructureType.buffer_image_copy2
	pNext             voidptr       = unsafe { nil }
	bufferOffset      DeviceSize
	bufferRowLength   u32
	bufferImageHeight u32
	imageSubresource  ImageSubresourceLayers
	imageOffset       Offset3D
	imageExtent       Extent3D
}

pub type CopyBufferToImageInfo2 = C.VkCopyBufferToImageInfo2

@[typedef]
pub struct C.VkCopyBufferToImageInfo2 {
pub mut:
	sType          StructureType = StructureType.copy_buffer_to_image_info2
	pNext          voidptr       = unsafe { nil }
	srcBuffer      Buffer
	dstImage       Image
	dstImageLayout ImageLayout
	regionCount    u32
	pRegions       &BufferImageCopy2
}

pub type CopyImageToBufferInfo2 = C.VkCopyImageToBufferInfo2

@[typedef]
pub struct C.VkCopyImageToBufferInfo2 {
pub mut:
	sType          StructureType = StructureType.copy_image_to_buffer_info2
	pNext          voidptr       = unsafe { nil }
	srcImage       Image
	srcImageLayout ImageLayout
	dstBuffer      Buffer
	regionCount    u32
	pRegions       &BufferImageCopy2
}

// PhysicalDeviceTextureCompressionASTCHDRFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceTextureCompressionASTCHDRFeatures = C.VkPhysicalDeviceTextureCompressionASTCHDRFeatures

@[typedef]
pub struct C.VkPhysicalDeviceTextureCompressionASTCHDRFeatures {
pub mut:
	sType                      StructureType = StructureType.physical_device_texture_compression_astc_hdr_features
	pNext                      voidptr       = unsafe { nil }
	textureCompressionASTC_HDR Bool32
}

// FormatProperties3 extends VkFormatProperties2
pub type FormatProperties3 = C.VkFormatProperties3

@[typedef]
pub struct C.VkFormatProperties3 {
pub mut:
	sType                 StructureType = StructureType.format_properties3
	pNext                 voidptr       = unsafe { nil }
	linearTilingFeatures  FormatFeatureFlags2
	optimalTilingFeatures FormatFeatureFlags2
	bufferFeatures        FormatFeatureFlags2
}

// PhysicalDeviceMaintenance4Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMaintenance4Features = C.VkPhysicalDeviceMaintenance4Features

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance4Features {
pub mut:
	sType        StructureType = StructureType.physical_device_maintenance4_features
	pNext        voidptr       = unsafe { nil }
	maintenance4 Bool32
}

// PhysicalDeviceMaintenance4Properties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMaintenance4Properties = C.VkPhysicalDeviceMaintenance4Properties

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance4Properties {
pub mut:
	sType         StructureType = StructureType.physical_device_maintenance4_properties
	pNext         voidptr       = unsafe { nil }
	maxBufferSize DeviceSize
}

pub type DeviceBufferMemoryRequirements = C.VkDeviceBufferMemoryRequirements

@[typedef]
pub struct C.VkDeviceBufferMemoryRequirements {
pub mut:
	sType       StructureType = StructureType.device_buffer_memory_requirements
	pNext       voidptr       = unsafe { nil }
	pCreateInfo &BufferCreateInfo
}

pub type DeviceImageMemoryRequirements = C.VkDeviceImageMemoryRequirements

@[typedef]
pub struct C.VkDeviceImageMemoryRequirements {
pub mut:
	sType       StructureType = StructureType.device_image_memory_requirements
	pNext       voidptr       = unsafe { nil }
	pCreateInfo &ImageCreateInfo
	planeAspect ImageAspectFlagBits
}

pub type PipelineCreationFeedback = C.VkPipelineCreationFeedback

@[typedef]
pub struct C.VkPipelineCreationFeedback {
pub mut:
	flags    PipelineCreationFeedbackFlags
	duration u64
}

// PipelineCreationFeedbackCreateInfo extends VkGraphicsPipelineCreateInfo,VkComputePipelineCreateInfo,VkRayTracingPipelineCreateInfoNV,VkRayTracingPipelineCreateInfoKHR,VkDataGraphPipelineCreateInfoARM
pub type PipelineCreationFeedbackCreateInfo = C.VkPipelineCreationFeedbackCreateInfo

@[typedef]
pub struct C.VkPipelineCreationFeedbackCreateInfo {
pub mut:
	sType                              StructureType = StructureType.pipeline_creation_feedback_create_info
	pNext                              voidptr       = unsafe { nil }
	pPipelineCreationFeedback          &PipelineCreationFeedback
	pipelineStageCreationFeedbackCount u32
	pPipelineStageCreationFeedbacks    &PipelineCreationFeedback
}

// PhysicalDeviceShaderTerminateInvocationFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderTerminateInvocationFeatures = C.VkPhysicalDeviceShaderTerminateInvocationFeatures

@[typedef]
pub struct C.VkPhysicalDeviceShaderTerminateInvocationFeatures {
pub mut:
	sType                     StructureType = StructureType.physical_device_shader_terminate_invocation_features
	pNext                     voidptr       = unsafe { nil }
	shaderTerminateInvocation Bool32
}

// PhysicalDeviceShaderDemoteToHelperInvocationFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderDemoteToHelperInvocationFeatures = C.VkPhysicalDeviceShaderDemoteToHelperInvocationFeatures

@[typedef]
pub struct C.VkPhysicalDeviceShaderDemoteToHelperInvocationFeatures {
pub mut:
	sType                          StructureType = StructureType.physical_device_shader_demote_to_helper_invocation_features
	pNext                          voidptr       = unsafe { nil }
	shaderDemoteToHelperInvocation Bool32
}

// PhysicalDevicePipelineCreationCacheControlFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePipelineCreationCacheControlFeatures = C.VkPhysicalDevicePipelineCreationCacheControlFeatures

@[typedef]
pub struct C.VkPhysicalDevicePipelineCreationCacheControlFeatures {
pub mut:
	sType                        StructureType = StructureType.physical_device_pipeline_creation_cache_control_features
	pNext                        voidptr       = unsafe { nil }
	pipelineCreationCacheControl Bool32
}

// PhysicalDeviceZeroInitializeWorkgroupMemoryFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceZeroInitializeWorkgroupMemoryFeatures = C.VkPhysicalDeviceZeroInitializeWorkgroupMemoryFeatures

@[typedef]
pub struct C.VkPhysicalDeviceZeroInitializeWorkgroupMemoryFeatures {
pub mut:
	sType                               StructureType = StructureType.physical_device_zero_initialize_workgroup_memory_features
	pNext                               voidptr       = unsafe { nil }
	shaderZeroInitializeWorkgroupMemory Bool32
}

// PhysicalDeviceImageRobustnessFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceImageRobustnessFeatures = C.VkPhysicalDeviceImageRobustnessFeatures

@[typedef]
pub struct C.VkPhysicalDeviceImageRobustnessFeatures {
pub mut:
	sType             StructureType = StructureType.physical_device_image_robustness_features
	pNext             voidptr       = unsafe { nil }
	robustImageAccess Bool32
}

// PhysicalDeviceSubgroupSizeControlFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceSubgroupSizeControlFeatures = C.VkPhysicalDeviceSubgroupSizeControlFeatures

@[typedef]
pub struct C.VkPhysicalDeviceSubgroupSizeControlFeatures {
pub mut:
	sType                StructureType = StructureType.physical_device_subgroup_size_control_features
	pNext                voidptr       = unsafe { nil }
	subgroupSizeControl  Bool32
	computeFullSubgroups Bool32
}

// PhysicalDeviceSubgroupSizeControlProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceSubgroupSizeControlProperties = C.VkPhysicalDeviceSubgroupSizeControlProperties

@[typedef]
pub struct C.VkPhysicalDeviceSubgroupSizeControlProperties {
pub mut:
	sType                        StructureType = StructureType.physical_device_subgroup_size_control_properties
	pNext                        voidptr       = unsafe { nil }
	minSubgroupSize              u32
	maxSubgroupSize              u32
	maxComputeWorkgroupSubgroups u32
	requiredSubgroupSizeStages   ShaderStageFlags
}

// PipelineShaderStageRequiredSubgroupSizeCreateInfo extends VkPipelineShaderStageCreateInfo,VkShaderCreateInfoEXT
pub type PipelineShaderStageRequiredSubgroupSizeCreateInfo = C.VkPipelineShaderStageRequiredSubgroupSizeCreateInfo

@[typedef]
pub struct C.VkPipelineShaderStageRequiredSubgroupSizeCreateInfo {
pub mut:
	sType                StructureType = StructureType.pipeline_shader_stage_required_subgroup_size_create_info
	pNext                voidptr       = unsafe { nil }
	requiredSubgroupSize u32
}

// PhysicalDeviceInlineUniformBlockFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceInlineUniformBlockFeatures = C.VkPhysicalDeviceInlineUniformBlockFeatures

@[typedef]
pub struct C.VkPhysicalDeviceInlineUniformBlockFeatures {
pub mut:
	sType                                              StructureType = StructureType.physical_device_inline_uniform_block_features
	pNext                                              voidptr       = unsafe { nil }
	inlineUniformBlock                                 Bool32
	descriptorBindingInlineUniformBlockUpdateAfterBind Bool32
}

// PhysicalDeviceInlineUniformBlockProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceInlineUniformBlockProperties = C.VkPhysicalDeviceInlineUniformBlockProperties

@[typedef]
pub struct C.VkPhysicalDeviceInlineUniformBlockProperties {
pub mut:
	sType                                                   StructureType = StructureType.physical_device_inline_uniform_block_properties
	pNext                                                   voidptr       = unsafe { nil }
	maxInlineUniformBlockSize                               u32
	maxPerStageDescriptorInlineUniformBlocks                u32
	maxPerStageDescriptorUpdateAfterBindInlineUniformBlocks u32
	maxDescriptorSetInlineUniformBlocks                     u32
	maxDescriptorSetUpdateAfterBindInlineUniformBlocks      u32
}

// WriteDescriptorSetInlineUniformBlock extends VkWriteDescriptorSet
pub type WriteDescriptorSetInlineUniformBlock = C.VkWriteDescriptorSetInlineUniformBlock

@[typedef]
pub struct C.VkWriteDescriptorSetInlineUniformBlock {
pub mut:
	sType    StructureType = StructureType.write_descriptor_set_inline_uniform_block
	pNext    voidptr       = unsafe { nil }
	dataSize u32
	pData    voidptr
}

// DescriptorPoolInlineUniformBlockCreateInfo extends VkDescriptorPoolCreateInfo
pub type DescriptorPoolInlineUniformBlockCreateInfo = C.VkDescriptorPoolInlineUniformBlockCreateInfo

@[typedef]
pub struct C.VkDescriptorPoolInlineUniformBlockCreateInfo {
pub mut:
	sType                         StructureType = StructureType.descriptor_pool_inline_uniform_block_create_info
	pNext                         voidptr       = unsafe { nil }
	maxInlineUniformBlockBindings u32
}

// PhysicalDeviceShaderIntegerDotProductFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderIntegerDotProductFeatures = C.VkPhysicalDeviceShaderIntegerDotProductFeatures

@[typedef]
pub struct C.VkPhysicalDeviceShaderIntegerDotProductFeatures {
pub mut:
	sType                   StructureType = StructureType.physical_device_shader_integer_dot_product_features
	pNext                   voidptr       = unsafe { nil }
	shaderIntegerDotProduct Bool32
}

// PhysicalDeviceShaderIntegerDotProductProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceShaderIntegerDotProductProperties = C.VkPhysicalDeviceShaderIntegerDotProductProperties

@[typedef]
pub struct C.VkPhysicalDeviceShaderIntegerDotProductProperties {
pub mut:
	sType                                                                         StructureType = StructureType.physical_device_shader_integer_dot_product_properties
	pNext                                                                         voidptr       = unsafe { nil }
	integerDotProduct8BitUnsignedAccelerated                                      Bool32
	integerDotProduct8BitSignedAccelerated                                        Bool32
	integerDotProduct8BitMixedSignednessAccelerated                               Bool32
	integerDotProduct4x8BitPackedUnsignedAccelerated                              Bool32
	integerDotProduct4x8BitPackedSignedAccelerated                                Bool32
	integerDotProduct4x8BitPackedMixedSignednessAccelerated                       Bool32
	integerDotProduct16BitUnsignedAccelerated                                     Bool32
	integerDotProduct16BitSignedAccelerated                                       Bool32
	integerDotProduct16BitMixedSignednessAccelerated                              Bool32
	integerDotProduct32BitUnsignedAccelerated                                     Bool32
	integerDotProduct32BitSignedAccelerated                                       Bool32
	integerDotProduct32BitMixedSignednessAccelerated                              Bool32
	integerDotProduct64BitUnsignedAccelerated                                     Bool32
	integerDotProduct64BitSignedAccelerated                                       Bool32
	integerDotProduct64BitMixedSignednessAccelerated                              Bool32
	integerDotProductAccumulatingSaturating8BitUnsignedAccelerated                Bool32
	integerDotProductAccumulatingSaturating8BitSignedAccelerated                  Bool32
	integerDotProductAccumulatingSaturating8BitMixedSignednessAccelerated         Bool32
	integerDotProductAccumulatingSaturating4x8BitPackedUnsignedAccelerated        Bool32
	integerDotProductAccumulatingSaturating4x8BitPackedSignedAccelerated          Bool32
	integerDotProductAccumulatingSaturating4x8BitPackedMixedSignednessAccelerated Bool32
	integerDotProductAccumulatingSaturating16BitUnsignedAccelerated               Bool32
	integerDotProductAccumulatingSaturating16BitSignedAccelerated                 Bool32
	integerDotProductAccumulatingSaturating16BitMixedSignednessAccelerated        Bool32
	integerDotProductAccumulatingSaturating32BitUnsignedAccelerated               Bool32
	integerDotProductAccumulatingSaturating32BitSignedAccelerated                 Bool32
	integerDotProductAccumulatingSaturating32BitMixedSignednessAccelerated        Bool32
	integerDotProductAccumulatingSaturating64BitUnsignedAccelerated               Bool32
	integerDotProductAccumulatingSaturating64BitSignedAccelerated                 Bool32
	integerDotProductAccumulatingSaturating64BitMixedSignednessAccelerated        Bool32
}

// PhysicalDeviceTexelBufferAlignmentProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceTexelBufferAlignmentProperties = C.VkPhysicalDeviceTexelBufferAlignmentProperties

@[typedef]
pub struct C.VkPhysicalDeviceTexelBufferAlignmentProperties {
pub mut:
	sType                                        StructureType = StructureType.physical_device_texel_buffer_alignment_properties
	pNext                                        voidptr       = unsafe { nil }
	storageTexelBufferOffsetAlignmentBytes       DeviceSize
	storageTexelBufferOffsetSingleTexelAlignment Bool32
	uniformTexelBufferOffsetAlignmentBytes       DeviceSize
	uniformTexelBufferOffsetSingleTexelAlignment Bool32
}

pub type ImageBlit2 = C.VkImageBlit2

@[typedef]
pub struct C.VkImageBlit2 {
pub mut:
	sType          StructureType = StructureType.image_blit2
	pNext          voidptr       = unsafe { nil }
	srcSubresource ImageSubresourceLayers
	srcOffsets     [2]Offset3D
	dstSubresource ImageSubresourceLayers
	dstOffsets     [2]Offset3D
}

pub type BlitImageInfo2 = C.VkBlitImageInfo2

@[typedef]
pub struct C.VkBlitImageInfo2 {
pub mut:
	sType          StructureType = StructureType.blit_image_info2
	pNext          voidptr       = unsafe { nil }
	srcImage       Image
	srcImageLayout ImageLayout
	dstImage       Image
	dstImageLayout ImageLayout
	regionCount    u32
	pRegions       &ImageBlit2
	filter         Filter
}

pub type ImageResolve2 = C.VkImageResolve2

@[typedef]
pub struct C.VkImageResolve2 {
pub mut:
	sType          StructureType = StructureType.image_resolve2
	pNext          voidptr       = unsafe { nil }
	srcSubresource ImageSubresourceLayers
	srcOffset      Offset3D
	dstSubresource ImageSubresourceLayers
	dstOffset      Offset3D
	extent         Extent3D
}

pub type ResolveImageInfo2 = C.VkResolveImageInfo2

@[typedef]
pub struct C.VkResolveImageInfo2 {
pub mut:
	sType          StructureType = StructureType.resolve_image_info2
	pNext          voidptr       = unsafe { nil }
	srcImage       Image
	srcImageLayout ImageLayout
	dstImage       Image
	dstImageLayout ImageLayout
	regionCount    u32
	pRegions       &ImageResolve2
}

pub type RenderingAttachmentInfo = C.VkRenderingAttachmentInfo

@[typedef]
pub struct C.VkRenderingAttachmentInfo {
pub mut:
	sType              StructureType = StructureType.rendering_attachment_info
	pNext              voidptr       = unsafe { nil }
	imageView          ImageView
	imageLayout        ImageLayout
	resolveMode        ResolveModeFlagBits
	resolveImageView   ImageView
	resolveImageLayout ImageLayout
	loadOp             AttachmentLoadOp
	storeOp            AttachmentStoreOp
	clearValue         ClearValue
}

pub type RenderingInfo = C.VkRenderingInfo

@[typedef]
pub struct C.VkRenderingInfo {
pub mut:
	sType                StructureType = StructureType.rendering_info
	pNext                voidptr       = unsafe { nil }
	flags                RenderingFlags
	renderArea           Rect2D
	layerCount           u32
	viewMask             u32
	colorAttachmentCount u32
	pColorAttachments    &RenderingAttachmentInfo
	pDepthAttachment     &RenderingAttachmentInfo
	pStencilAttachment   &RenderingAttachmentInfo
}

// PipelineRenderingCreateInfo extends VkGraphicsPipelineCreateInfo
pub type PipelineRenderingCreateInfo = C.VkPipelineRenderingCreateInfo

@[typedef]
pub struct C.VkPipelineRenderingCreateInfo {
pub mut:
	sType                   StructureType = StructureType.pipeline_rendering_create_info
	pNext                   voidptr       = unsafe { nil }
	viewMask                u32
	colorAttachmentCount    u32
	pColorAttachmentFormats &Format
	depthAttachmentFormat   Format
	stencilAttachmentFormat Format
}

// PhysicalDeviceDynamicRenderingFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDynamicRenderingFeatures = C.VkPhysicalDeviceDynamicRenderingFeatures

@[typedef]
pub struct C.VkPhysicalDeviceDynamicRenderingFeatures {
pub mut:
	sType            StructureType = StructureType.physical_device_dynamic_rendering_features
	pNext            voidptr       = unsafe { nil }
	dynamicRendering Bool32
}

// CommandBufferInheritanceRenderingInfo extends VkCommandBufferInheritanceInfo
pub type CommandBufferInheritanceRenderingInfo = C.VkCommandBufferInheritanceRenderingInfo

@[typedef]
pub struct C.VkCommandBufferInheritanceRenderingInfo {
pub mut:
	sType                   StructureType = StructureType.command_buffer_inheritance_rendering_info
	pNext                   voidptr       = unsafe { nil }
	flags                   RenderingFlags
	viewMask                u32
	colorAttachmentCount    u32
	pColorAttachmentFormats &Format
	depthAttachmentFormat   Format
	stencilAttachmentFormat Format
	rasterizationSamples    SampleCountFlagBits
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceToolProperties(physical_device PhysicalDevice, p_tool_count &u32, mut p_tool_properties PhysicalDeviceToolProperties) Result

pub type PFN_vkGetPhysicalDeviceToolProperties = fn (physical_device PhysicalDevice, p_tool_count &u32, mut p_tool_properties PhysicalDeviceToolProperties) Result

@[inline]
pub fn get_physical_device_tool_properties(physical_device PhysicalDevice,
	p_tool_count &u32,
	mut p_tool_properties PhysicalDeviceToolProperties) Result {
	return C.vkGetPhysicalDeviceToolProperties(physical_device, p_tool_count, mut p_tool_properties)
}

@[keep_args_alive]
fn C.vkCreatePrivateDataSlot(device Device, p_create_info &PrivateDataSlotCreateInfo, p_allocator &AllocationCallbacks, p_private_data_slot &PrivateDataSlot) Result

pub type PFN_vkCreatePrivateDataSlot = fn (device Device, p_create_info &PrivateDataSlotCreateInfo, p_allocator &AllocationCallbacks, p_private_data_slot &PrivateDataSlot) Result

@[inline]
pub fn create_private_data_slot(device Device,
	p_create_info &PrivateDataSlotCreateInfo,
	p_allocator &AllocationCallbacks,
	p_private_data_slot &PrivateDataSlot) Result {
	return C.vkCreatePrivateDataSlot(device, p_create_info, p_allocator, p_private_data_slot)
}

@[keep_args_alive]
fn C.vkDestroyPrivateDataSlot(device Device, private_data_slot PrivateDataSlot, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyPrivateDataSlot = fn (device Device, private_data_slot PrivateDataSlot, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_private_data_slot(device Device,
	private_data_slot PrivateDataSlot,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyPrivateDataSlot(device, private_data_slot, p_allocator)
}

@[keep_args_alive]
fn C.vkSetPrivateData(device Device, object_type ObjectType, object_handle u64, private_data_slot PrivateDataSlot, data u64) Result

pub type PFN_vkSetPrivateData = fn (device Device, object_type ObjectType, object_handle u64, private_data_slot PrivateDataSlot, data u64) Result

@[inline]
pub fn set_private_data(device Device,
	object_type ObjectType,
	object_handle u64,
	private_data_slot PrivateDataSlot,
	data u64) Result {
	return C.vkSetPrivateData(device, object_type, object_handle, private_data_slot, data)
}

@[keep_args_alive]
fn C.vkGetPrivateData(device Device, object_type ObjectType, object_handle u64, private_data_slot PrivateDataSlot, p_data &u64)

pub type PFN_vkGetPrivateData = fn (device Device, object_type ObjectType, object_handle u64, private_data_slot PrivateDataSlot, p_data &u64)

@[inline]
pub fn get_private_data(device Device,
	object_type ObjectType,
	object_handle u64,
	private_data_slot PrivateDataSlot,
	p_data &u64) {
	C.vkGetPrivateData(device, object_type, object_handle, private_data_slot, p_data)
}

@[keep_args_alive]
fn C.vkCmdPipelineBarrier2(command_buffer CommandBuffer, p_dependency_info &DependencyInfo)

pub type PFN_vkCmdPipelineBarrier2 = fn (command_buffer CommandBuffer, p_dependency_info &DependencyInfo)

@[inline]
pub fn cmd_pipeline_barrier2(command_buffer CommandBuffer,
	p_dependency_info &DependencyInfo) {
	C.vkCmdPipelineBarrier2(command_buffer, p_dependency_info)
}

@[keep_args_alive]
fn C.vkCmdWriteTimestamp2(command_buffer CommandBuffer, stage PipelineStageFlags2, query_pool QueryPool, query u32)

pub type PFN_vkCmdWriteTimestamp2 = fn (command_buffer CommandBuffer, stage PipelineStageFlags2, query_pool QueryPool, query u32)

@[inline]
pub fn cmd_write_timestamp2(command_buffer CommandBuffer,
	stage PipelineStageFlags2,
	query_pool QueryPool,
	query u32) {
	C.vkCmdWriteTimestamp2(command_buffer, stage, query_pool, query)
}

@[keep_args_alive]
fn C.vkQueueSubmit2(queue Queue, submit_count u32, p_submits &SubmitInfo2, fence Fence) Result

pub type PFN_vkQueueSubmit2 = fn (queue Queue, submit_count u32, p_submits &SubmitInfo2, fence Fence) Result

@[inline]
pub fn queue_submit2(queue Queue,
	submit_count u32,
	p_submits &SubmitInfo2,
	fence Fence) Result {
	return C.vkQueueSubmit2(queue, submit_count, p_submits, fence)
}

@[keep_args_alive]
fn C.vkCmdCopyBuffer2(command_buffer CommandBuffer, p_copy_buffer_info &CopyBufferInfo2)

pub type PFN_vkCmdCopyBuffer2 = fn (command_buffer CommandBuffer, p_copy_buffer_info &CopyBufferInfo2)

@[inline]
pub fn cmd_copy_buffer2(command_buffer CommandBuffer,
	p_copy_buffer_info &CopyBufferInfo2) {
	C.vkCmdCopyBuffer2(command_buffer, p_copy_buffer_info)
}

@[keep_args_alive]
fn C.vkCmdCopyImage2(command_buffer CommandBuffer, p_copy_image_info &CopyImageInfo2)

pub type PFN_vkCmdCopyImage2 = fn (command_buffer CommandBuffer, p_copy_image_info &CopyImageInfo2)

@[inline]
pub fn cmd_copy_image2(command_buffer CommandBuffer,
	p_copy_image_info &CopyImageInfo2) {
	C.vkCmdCopyImage2(command_buffer, p_copy_image_info)
}

@[keep_args_alive]
fn C.vkCmdCopyBufferToImage2(command_buffer CommandBuffer, p_copy_buffer_to_image_info &CopyBufferToImageInfo2)

pub type PFN_vkCmdCopyBufferToImage2 = fn (command_buffer CommandBuffer, p_copy_buffer_to_image_info &CopyBufferToImageInfo2)

@[inline]
pub fn cmd_copy_buffer_to_image2(command_buffer CommandBuffer,
	p_copy_buffer_to_image_info &CopyBufferToImageInfo2) {
	C.vkCmdCopyBufferToImage2(command_buffer, p_copy_buffer_to_image_info)
}

@[keep_args_alive]
fn C.vkCmdCopyImageToBuffer2(command_buffer CommandBuffer, p_copy_image_to_buffer_info &CopyImageToBufferInfo2)

pub type PFN_vkCmdCopyImageToBuffer2 = fn (command_buffer CommandBuffer, p_copy_image_to_buffer_info &CopyImageToBufferInfo2)

@[inline]
pub fn cmd_copy_image_to_buffer2(command_buffer CommandBuffer,
	p_copy_image_to_buffer_info &CopyImageToBufferInfo2) {
	C.vkCmdCopyImageToBuffer2(command_buffer, p_copy_image_to_buffer_info)
}

@[keep_args_alive]
fn C.vkGetDeviceBufferMemoryRequirements(device Device, p_info &DeviceBufferMemoryRequirements, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetDeviceBufferMemoryRequirements = fn (device Device, p_info &DeviceBufferMemoryRequirements, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_device_buffer_memory_requirements(device Device,
	p_info &DeviceBufferMemoryRequirements,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetDeviceBufferMemoryRequirements(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetDeviceImageMemoryRequirements(device Device, p_info &DeviceImageMemoryRequirements, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetDeviceImageMemoryRequirements = fn (device Device, p_info &DeviceImageMemoryRequirements, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_device_image_memory_requirements(device Device,
	p_info &DeviceImageMemoryRequirements,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetDeviceImageMemoryRequirements(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetDeviceImageSparseMemoryRequirements(device Device, p_info &DeviceImageMemoryRequirements, p_sparse_memory_requirement_count &u32, mut p_sparse_memory_requirements SparseImageMemoryRequirements2)

pub type PFN_vkGetDeviceImageSparseMemoryRequirements = fn (device Device, p_info &DeviceImageMemoryRequirements, p_sparse_memory_requirement_count &u32, mut p_sparse_memory_requirements SparseImageMemoryRequirements2)

@[inline]
pub fn get_device_image_sparse_memory_requirements(device Device,
	p_info &DeviceImageMemoryRequirements,
	p_sparse_memory_requirement_count &u32,
	mut p_sparse_memory_requirements SparseImageMemoryRequirements2) {
	C.vkGetDeviceImageSparseMemoryRequirements(device, p_info, p_sparse_memory_requirement_count, mut
		p_sparse_memory_requirements)
}

@[keep_args_alive]
fn C.vkCmdSetEvent2(command_buffer CommandBuffer, event Event, p_dependency_info &DependencyInfo)

pub type PFN_vkCmdSetEvent2 = fn (command_buffer CommandBuffer, event Event, p_dependency_info &DependencyInfo)

@[inline]
pub fn cmd_set_event2(command_buffer CommandBuffer,
	event Event,
	p_dependency_info &DependencyInfo) {
	C.vkCmdSetEvent2(command_buffer, event, p_dependency_info)
}

@[keep_args_alive]
fn C.vkCmdResetEvent2(command_buffer CommandBuffer, event Event, stage_mask PipelineStageFlags2)

pub type PFN_vkCmdResetEvent2 = fn (command_buffer CommandBuffer, event Event, stage_mask PipelineStageFlags2)

@[inline]
pub fn cmd_reset_event2(command_buffer CommandBuffer,
	event Event,
	stage_mask PipelineStageFlags2) {
	C.vkCmdResetEvent2(command_buffer, event, stage_mask)
}

@[keep_args_alive]
fn C.vkCmdWaitEvents2(command_buffer CommandBuffer, event_count u32, p_events &Event, p_dependency_infos &DependencyInfo)

pub type PFN_vkCmdWaitEvents2 = fn (command_buffer CommandBuffer, event_count u32, p_events &Event, p_dependency_infos &DependencyInfo)

@[inline]
pub fn cmd_wait_events2(command_buffer CommandBuffer,
	event_count u32,
	p_events &Event,
	p_dependency_infos &DependencyInfo) {
	C.vkCmdWaitEvents2(command_buffer, event_count, p_events, p_dependency_infos)
}

@[keep_args_alive]
fn C.vkCmdBlitImage2(command_buffer CommandBuffer, p_blit_image_info &BlitImageInfo2)

pub type PFN_vkCmdBlitImage2 = fn (command_buffer CommandBuffer, p_blit_image_info &BlitImageInfo2)

@[inline]
pub fn cmd_blit_image2(command_buffer CommandBuffer,
	p_blit_image_info &BlitImageInfo2) {
	C.vkCmdBlitImage2(command_buffer, p_blit_image_info)
}

@[keep_args_alive]
fn C.vkCmdResolveImage2(command_buffer CommandBuffer, p_resolve_image_info &ResolveImageInfo2)

pub type PFN_vkCmdResolveImage2 = fn (command_buffer CommandBuffer, p_resolve_image_info &ResolveImageInfo2)

@[inline]
pub fn cmd_resolve_image2(command_buffer CommandBuffer,
	p_resolve_image_info &ResolveImageInfo2) {
	C.vkCmdResolveImage2(command_buffer, p_resolve_image_info)
}

@[keep_args_alive]
fn C.vkCmdBeginRendering(command_buffer CommandBuffer, p_rendering_info &RenderingInfo)

pub type PFN_vkCmdBeginRendering = fn (command_buffer CommandBuffer, p_rendering_info &RenderingInfo)

@[inline]
pub fn cmd_begin_rendering(command_buffer CommandBuffer,
	p_rendering_info &RenderingInfo) {
	C.vkCmdBeginRendering(command_buffer, p_rendering_info)
}

@[keep_args_alive]
fn C.vkCmdEndRendering(command_buffer CommandBuffer)

pub type PFN_vkCmdEndRendering = fn (command_buffer CommandBuffer)

@[inline]
pub fn cmd_end_rendering(command_buffer CommandBuffer) {
	C.vkCmdEndRendering(command_buffer)
}

@[keep_args_alive]
fn C.vkCmdSetCullMode(command_buffer CommandBuffer, cull_mode CullModeFlags)

pub type PFN_vkCmdSetCullMode = fn (command_buffer CommandBuffer, cull_mode CullModeFlags)

@[inline]
pub fn cmd_set_cull_mode(command_buffer CommandBuffer,
	cull_mode CullModeFlags) {
	C.vkCmdSetCullMode(command_buffer, cull_mode)
}

@[keep_args_alive]
fn C.vkCmdSetFrontFace(command_buffer CommandBuffer, front_face FrontFace)

pub type PFN_vkCmdSetFrontFace = fn (command_buffer CommandBuffer, front_face FrontFace)

@[inline]
pub fn cmd_set_front_face(command_buffer CommandBuffer,
	front_face FrontFace) {
	C.vkCmdSetFrontFace(command_buffer, front_face)
}

@[keep_args_alive]
fn C.vkCmdSetPrimitiveTopology(command_buffer CommandBuffer, primitive_topology PrimitiveTopology)

pub type PFN_vkCmdSetPrimitiveTopology = fn (command_buffer CommandBuffer, primitive_topology PrimitiveTopology)

@[inline]
pub fn cmd_set_primitive_topology(command_buffer CommandBuffer,
	primitive_topology PrimitiveTopology) {
	C.vkCmdSetPrimitiveTopology(command_buffer, primitive_topology)
}

@[keep_args_alive]
fn C.vkCmdSetViewportWithCount(command_buffer CommandBuffer, viewport_count u32, p_viewports &Viewport)

pub type PFN_vkCmdSetViewportWithCount = fn (command_buffer CommandBuffer, viewport_count u32, p_viewports &Viewport)

@[inline]
pub fn cmd_set_viewport_with_count(command_buffer CommandBuffer,
	viewport_count u32,
	p_viewports &Viewport) {
	C.vkCmdSetViewportWithCount(command_buffer, viewport_count, p_viewports)
}

@[keep_args_alive]
fn C.vkCmdSetScissorWithCount(command_buffer CommandBuffer, scissor_count u32, p_scissors &Rect2D)

pub type PFN_vkCmdSetScissorWithCount = fn (command_buffer CommandBuffer, scissor_count u32, p_scissors &Rect2D)

@[inline]
pub fn cmd_set_scissor_with_count(command_buffer CommandBuffer,
	scissor_count u32,
	p_scissors &Rect2D) {
	C.vkCmdSetScissorWithCount(command_buffer, scissor_count, p_scissors)
}

@[keep_args_alive]
fn C.vkCmdBindVertexBuffers2(command_buffer CommandBuffer, first_binding u32, binding_count u32, p_buffers &Buffer, p_offsets &DeviceSize, p_sizes &DeviceSize, p_strides &DeviceSize)

pub type PFN_vkCmdBindVertexBuffers2 = fn (command_buffer CommandBuffer, first_binding u32, binding_count u32, p_buffers &Buffer, p_offsets &DeviceSize, p_sizes &DeviceSize, p_strides &DeviceSize)

@[inline]
pub fn cmd_bind_vertex_buffers2(command_buffer CommandBuffer,
	first_binding u32,
	binding_count u32,
	p_buffers &Buffer,
	p_offsets &DeviceSize,
	p_sizes &DeviceSize,
	p_strides &DeviceSize) {
	C.vkCmdBindVertexBuffers2(command_buffer, first_binding, binding_count, p_buffers,
		p_offsets, p_sizes, p_strides)
}

@[keep_args_alive]
fn C.vkCmdSetDepthTestEnable(command_buffer CommandBuffer, depth_test_enable Bool32)

pub type PFN_vkCmdSetDepthTestEnable = fn (command_buffer CommandBuffer, depth_test_enable Bool32)

@[inline]
pub fn cmd_set_depth_test_enable(command_buffer CommandBuffer,
	depth_test_enable Bool32) {
	C.vkCmdSetDepthTestEnable(command_buffer, depth_test_enable)
}

@[keep_args_alive]
fn C.vkCmdSetDepthWriteEnable(command_buffer CommandBuffer, depth_write_enable Bool32)

pub type PFN_vkCmdSetDepthWriteEnable = fn (command_buffer CommandBuffer, depth_write_enable Bool32)

@[inline]
pub fn cmd_set_depth_write_enable(command_buffer CommandBuffer,
	depth_write_enable Bool32) {
	C.vkCmdSetDepthWriteEnable(command_buffer, depth_write_enable)
}

@[keep_args_alive]
fn C.vkCmdSetDepthCompareOp(command_buffer CommandBuffer, depth_compare_op CompareOp)

pub type PFN_vkCmdSetDepthCompareOp = fn (command_buffer CommandBuffer, depth_compare_op CompareOp)

@[inline]
pub fn cmd_set_depth_compare_op(command_buffer CommandBuffer,
	depth_compare_op CompareOp) {
	C.vkCmdSetDepthCompareOp(command_buffer, depth_compare_op)
}

@[keep_args_alive]
fn C.vkCmdSetDepthBoundsTestEnable(command_buffer CommandBuffer, depth_bounds_test_enable Bool32)

pub type PFN_vkCmdSetDepthBoundsTestEnable = fn (command_buffer CommandBuffer, depth_bounds_test_enable Bool32)

@[inline]
pub fn cmd_set_depth_bounds_test_enable(command_buffer CommandBuffer,
	depth_bounds_test_enable Bool32) {
	C.vkCmdSetDepthBoundsTestEnable(command_buffer, depth_bounds_test_enable)
}

@[keep_args_alive]
fn C.vkCmdSetStencilTestEnable(command_buffer CommandBuffer, stencil_test_enable Bool32)

pub type PFN_vkCmdSetStencilTestEnable = fn (command_buffer CommandBuffer, stencil_test_enable Bool32)

@[inline]
pub fn cmd_set_stencil_test_enable(command_buffer CommandBuffer,
	stencil_test_enable Bool32) {
	C.vkCmdSetStencilTestEnable(command_buffer, stencil_test_enable)
}

@[keep_args_alive]
fn C.vkCmdSetStencilOp(command_buffer CommandBuffer, face_mask StencilFaceFlags, fail_op StencilOp, pass_op StencilOp, depth_fail_op StencilOp, compare_op CompareOp)

pub type PFN_vkCmdSetStencilOp = fn (command_buffer CommandBuffer, face_mask StencilFaceFlags, fail_op StencilOp, pass_op StencilOp, depth_fail_op StencilOp, compare_op CompareOp)

@[inline]
pub fn cmd_set_stencil_op(command_buffer CommandBuffer,
	face_mask StencilFaceFlags,
	fail_op StencilOp,
	pass_op StencilOp,
	depth_fail_op StencilOp,
	compare_op CompareOp) {
	C.vkCmdSetStencilOp(command_buffer, face_mask, fail_op, pass_op, depth_fail_op, compare_op)
}

@[keep_args_alive]
fn C.vkCmdSetRasterizerDiscardEnable(command_buffer CommandBuffer, rasterizer_discard_enable Bool32)

pub type PFN_vkCmdSetRasterizerDiscardEnable = fn (command_buffer CommandBuffer, rasterizer_discard_enable Bool32)

@[inline]
pub fn cmd_set_rasterizer_discard_enable(command_buffer CommandBuffer,
	rasterizer_discard_enable Bool32) {
	C.vkCmdSetRasterizerDiscardEnable(command_buffer, rasterizer_discard_enable)
}

@[keep_args_alive]
fn C.vkCmdSetDepthBiasEnable(command_buffer CommandBuffer, depth_bias_enable Bool32)

pub type PFN_vkCmdSetDepthBiasEnable = fn (command_buffer CommandBuffer, depth_bias_enable Bool32)

@[inline]
pub fn cmd_set_depth_bias_enable(command_buffer CommandBuffer,
	depth_bias_enable Bool32) {
	C.vkCmdSetDepthBiasEnable(command_buffer, depth_bias_enable)
}

@[keep_args_alive]
fn C.vkCmdSetPrimitiveRestartEnable(command_buffer CommandBuffer, primitive_restart_enable Bool32)

pub type PFN_vkCmdSetPrimitiveRestartEnable = fn (command_buffer CommandBuffer, primitive_restart_enable Bool32)

@[inline]
pub fn cmd_set_primitive_restart_enable(command_buffer CommandBuffer,
	primitive_restart_enable Bool32) {
	C.vkCmdSetPrimitiveRestartEnable(command_buffer, primitive_restart_enable)
}

pub const api_version_1_4 = make_api_version(0, 1, 4, 0) // patch version should always be set to 0
pub const max_global_priority_size = u32(16)

pub enum PipelineRobustnessBufferBehavior as u32 {
	device_default        = 0
	disabled              = 1
	robust_buffer_access  = 2
	robust_buffer_access2 = 3
	max_enum              = max_int
}

pub enum PipelineRobustnessImageBehavior as u32 {
	device_default       = 0
	disabled             = 1
	robust_image_access  = 2
	robust_image_access2 = 3
	max_enum             = max_int
}

pub enum QueueGlobalPriority as u32 {
	low      = 128
	medium   = 256
	high     = 512
	realtime = 1024
	max_enum = max_int
}

pub enum LineRasterizationMode as u32 {
	default            = 0
	rectangular        = 1
	bresenham          = 2
	rectangular_smooth = 3
	max_enum           = max_int
}

pub enum MemoryUnmapFlagBits as u32 {
	reserve_bit_ext = u32(0x00000001)
	max_enum        = max_int
}
pub type MemoryUnmapFlags = u32
pub type BufferUsageFlags2 = u64

// Flag bits for BufferUsageFlagBits2
pub type BufferUsageFlagBits2 = u64

pub const buffer_usage_2_transfer_src_bit = u64(0x00000001)
pub const buffer_usage_2_transfer_dst_bit = u64(0x00000002)
pub const buffer_usage_2_uniform_texel_buffer_bit = u64(0x00000004)
pub const buffer_usage_2_storage_texel_buffer_bit = u64(0x00000008)
pub const buffer_usage_2_uniform_buffer_bit = u64(0x00000010)
pub const buffer_usage_2_storage_buffer_bit = u64(0x00000020)
pub const buffer_usage_2_index_buffer_bit = u64(0x00000040)
pub const buffer_usage_2_vertex_buffer_bit = u64(0x00000080)
pub const buffer_usage_2_indirect_buffer_bit = u64(0x00000100)
pub const buffer_usage_2_shader_device_address_bit = u64(0x00020000)
pub const buffer_usage_2_execution_graph_scratch_bit_amdx = u64(0x02000000)
pub const buffer_usage_2_transfer_src_bit_khr = u32(buffer_usage_2_transfer_src_bit)
pub const buffer_usage_2_transfer_dst_bit_khr = u32(buffer_usage_2_transfer_dst_bit)
pub const buffer_usage_2_uniform_texel_buffer_bit_khr = u32(buffer_usage_2_uniform_texel_buffer_bit)
pub const buffer_usage_2_storage_texel_buffer_bit_khr = u32(buffer_usage_2_storage_texel_buffer_bit)
pub const buffer_usage_2_uniform_buffer_bit_khr = u32(buffer_usage_2_uniform_buffer_bit)
pub const buffer_usage_2_storage_buffer_bit_khr = u32(buffer_usage_2_storage_buffer_bit)
pub const buffer_usage_2_index_buffer_bit_khr = u32(buffer_usage_2_index_buffer_bit)
pub const buffer_usage_2_vertex_buffer_bit_khr = u32(buffer_usage_2_vertex_buffer_bit)
pub const buffer_usage_2_indirect_buffer_bit_khr = u32(buffer_usage_2_indirect_buffer_bit)
pub const buffer_usage_2_conditional_rendering_bit_ext = u64(0x00000200)
pub const buffer_usage_2_shader_binding_table_bit_khr = u64(0x00000400)
pub const buffer_usage_2_ray_tracing_bit_nv = u32(buffer_usage_2_shader_binding_table_bit_khr)
pub const buffer_usage_2_transform_feedback_buffer_bit_ext = u64(0x00000800)
pub const buffer_usage_2_transform_feedback_counter_buffer_bit_ext = u64(0x00001000)
pub const buffer_usage_2_video_decode_src_bit_khr = u64(0x00002000)
pub const buffer_usage_2_video_decode_dst_bit_khr = u64(0x00004000)
pub const buffer_usage_2_video_encode_dst_bit_khr = u64(0x00008000)
pub const buffer_usage_2_video_encode_src_bit_khr = u64(0x00010000)
pub const buffer_usage_2_shader_device_address_bit_khr = u32(buffer_usage_2_shader_device_address_bit)
pub const buffer_usage_2_acceleration_structure_build_input_read_only_bit_khr = u64(0x00080000)
pub const buffer_usage_2_acceleration_structure_storage_bit_khr = u64(0x00100000)
pub const buffer_usage_2_sampler_descriptor_buffer_bit_ext = u64(0x00200000)
pub const buffer_usage_2_resource_descriptor_buffer_bit_ext = u64(0x00400000)
pub const buffer_usage_2_push_descriptors_descriptor_buffer_bit_ext = u64(0x04000000)
pub const buffer_usage_2_micromap_build_input_read_only_bit_ext = u64(0x00800000)
pub const buffer_usage_2_micromap_storage_bit_ext = u64(0x01000000)
pub const buffer_usage_2_compressed_data_dgf1_bit_amdx = u64(0x200000000)
pub const buffer_usage_2_data_graph_foreign_descriptor_bit_arm = u64(0x20000000)
pub const buffer_usage_2_tile_memory_bit_qcom = u64(0x08000000)
pub const buffer_usage_2_memory_decompression_bit_ext = u64(0x100000000)
pub const buffer_usage_2_preprocess_buffer_bit_ext = u64(0x80000000)

pub enum HostImageCopyFlagBits as u32 {
	memcpy   = u32(0x00000001)
	max_enum = max_int
}
pub type HostImageCopyFlags = u32
pub type PipelineCreateFlags2 = u64

// Flag bits for PipelineCreateFlagBits2
pub type PipelineCreateFlagBits2 = u64

pub const pipeline_create_2_disable_optimization_bit = u64(0x00000001)
pub const pipeline_create_2_allow_derivatives_bit = u64(0x00000002)
pub const pipeline_create_2_derivative_bit = u64(0x00000004)
pub const pipeline_create_2_view_index_from_device_index_bit = u64(0x00000008)
pub const pipeline_create_2_dispatch_base_bit = u64(0x00000010)
pub const pipeline_create_2_fail_on_pipeline_compile_required_bit = u64(0x00000100)
pub const pipeline_create_2_early_return_on_failure_bit = u64(0x00000200)
pub const pipeline_create_2_no_protected_access_bit = u64(0x08000000)
pub const pipeline_create_2_protected_access_only_bit = u64(0x40000000)
pub const pipeline_create_2_execution_graph_bit_amdx = u64(0x100000000)
pub const pipeline_create_2_ray_tracing_skip_built_in_primitives_bit_khr = pipeline_create_2_ray_tracing_skip_triangles_bit_khr
pub const pipeline_create_2_ray_tracing_allow_spheres_and_linear_swept_spheres_bit_nv = u64(0x200000000)
pub const pipeline_create_2_enable_legacy_dithering_bit_ext = u64(0x400000000)
pub const pipeline_create_2_disable_optimization_bit_khr = pipeline_create_2_disable_optimization_bit
pub const pipeline_create_2_allow_derivatives_bit_khr = pipeline_create_2_allow_derivatives_bit
pub const pipeline_create_2_derivative_bit_khr = pipeline_create_2_derivative_bit
pub const pipeline_create_2_view_index_from_device_index_bit_khr = pipeline_create_2_view_index_from_device_index_bit
pub const pipeline_create_2_dispatch_base_bit_khr = pipeline_create_2_dispatch_base_bit
pub const pipeline_create_2_defer_compile_bit_nv = u64(0x00000020)
pub const pipeline_create_2_capture_statistics_bit_khr = u64(0x00000040)
pub const pipeline_create_2_capture_internal_representations_bit_khr = u64(0x00000080)
pub const pipeline_create_2_fail_on_pipeline_compile_required_bit_khr = u32(pipeline_create_2_fail_on_pipeline_compile_required_bit)
pub const pipeline_create_2_early_return_on_failure_bit_khr = u32(pipeline_create_2_early_return_on_failure_bit)
pub const pipeline_create_2_link_time_optimization_bit_ext = u64(0x00000400)
pub const pipeline_create_2_retain_link_time_optimization_info_bit_ext = u64(0x00800000)
pub const pipeline_create_2_library_bit_khr = u64(0x00000800)
pub const pipeline_create_2_ray_tracing_skip_triangles_bit_khr = u64(0x00001000)
pub const pipeline_create_2_ray_tracing_skip_aabbs_bit_khr = u64(0x00002000)
pub const pipeline_create_2_ray_tracing_no_null_any_hit_shaders_bit_khr = u64(0x00004000)
pub const pipeline_create_2_ray_tracing_no_null_closest_hit_shaders_bit_khr = u64(0x00008000)
pub const pipeline_create_2_ray_tracing_no_null_miss_shaders_bit_khr = u64(0x00010000)
pub const pipeline_create_2_ray_tracing_no_null_intersection_shaders_bit_khr = u64(0x00020000)
pub const pipeline_create_2_ray_tracing_shader_group_handle_capture_replay_bit_khr = u64(0x00080000)
pub const pipeline_create_2_indirect_bindable_bit_nv = u64(0x00040000)
pub const pipeline_create_2_ray_tracing_allow_motion_bit_nv = u64(0x00100000)
pub const pipeline_create_2_rendering_fragment_shading_rate_attachment_bit_khr = u64(0x00200000)
pub const pipeline_create_2_rendering_fragment_density_map_attachment_bit_ext = u64(0x00400000)
pub const pipeline_create_2_ray_tracing_opacity_micromap_bit_ext = u64(0x01000000)
pub const pipeline_create_2_color_attachment_feedback_loop_bit_ext = u64(0x02000000)
pub const pipeline_create_2_depth_stencil_attachment_feedback_loop_bit_ext = u64(0x04000000)
pub const pipeline_create_2_no_protected_access_bit_ext = pipeline_create_2_no_protected_access_bit
pub const pipeline_create_2_protected_access_only_bit_ext = pipeline_create_2_protected_access_only_bit
pub const pipeline_create_2_ray_tracing_displacement_micromap_bit_nv = u64(0x10000000)
pub const pipeline_create_2_descriptor_buffer_bit_ext = u64(0x20000000)
pub const pipeline_create_2_disallow_opacity_micromap_bit_arm = u64(0x2000000000)
pub const pipeline_create_2_capture_data_bit_khr = u64(0x80000000)
pub const pipeline_create_2_indirect_bindable_bit_ext = u64(0x4000000000)
pub const pipeline_create_2_per_layer_fragment_density_bit_valve = u64(0x10000000000)
pub const pipeline_create_2_64_bit_indexing_bit_ext = u64(0x80000000000)

// PhysicalDeviceVulkan14Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVulkan14Features = C.VkPhysicalDeviceVulkan14Features

@[typedef]
pub struct C.VkPhysicalDeviceVulkan14Features {
pub mut:
	sType                                  StructureType = StructureType.physical_device_vulkan1_4_features
	pNext                                  voidptr       = unsafe { nil }
	globalPriorityQuery                    Bool32
	shaderSubgroupRotate                   Bool32
	shaderSubgroupRotateClustered          Bool32
	shaderFloatControls2                   Bool32
	shaderExpectAssume                     Bool32
	rectangularLines                       Bool32
	bresenhamLines                         Bool32
	smoothLines                            Bool32
	stippledRectangularLines               Bool32
	stippledBresenhamLines                 Bool32
	stippledSmoothLines                    Bool32
	vertexAttributeInstanceRateDivisor     Bool32
	vertexAttributeInstanceRateZeroDivisor Bool32
	indexTypeUint8                         Bool32
	dynamicRenderingLocalRead              Bool32
	maintenance5                           Bool32
	maintenance6                           Bool32
	pipelineProtectedAccess                Bool32
	pipelineRobustness                     Bool32
	hostImageCopy                          Bool32
	pushDescriptor                         Bool32
}

// PhysicalDeviceVulkan14Properties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceVulkan14Properties = C.VkPhysicalDeviceVulkan14Properties

@[typedef]
pub struct C.VkPhysicalDeviceVulkan14Properties {
pub mut:
	sType                                               StructureType = StructureType.physical_device_vulkan1_4_properties
	pNext                                               voidptr       = unsafe { nil }
	lineSubPixelPrecisionBits                           u32
	maxVertexAttribDivisor                              u32
	supportsNonZeroFirstInstance                        Bool32
	maxPushDescriptors                                  u32
	dynamicRenderingLocalReadDepthStencilAttachments    Bool32
	dynamicRenderingLocalReadMultisampledAttachments    Bool32
	earlyFragmentMultisampleCoverageAfterSampleCounting Bool32
	earlyFragmentSampleMaskTestBeforeSampleCounting     Bool32
	depthStencilSwizzleOneSupport                       Bool32
	polygonModePointSize                                Bool32
	nonStrictSinglePixelWideLinesUseParallelogram       Bool32
	nonStrictWideLinesUseParallelogram                  Bool32
	blockTexelViewCompatibleMultipleLayers              Bool32
	maxCombinedImageSamplerDescriptorCount              u32
	fragmentShadingRateClampCombinerInputs              Bool32
	defaultRobustnessStorageBuffers                     PipelineRobustnessBufferBehavior
	defaultRobustnessUniformBuffers                     PipelineRobustnessBufferBehavior
	defaultRobustnessVertexInputs                       PipelineRobustnessBufferBehavior
	defaultRobustnessImages                             PipelineRobustnessImageBehavior
	copySrcLayoutCount                                  u32
	pCopySrcLayouts                                     &ImageLayout
	copyDstLayoutCount                                  u32
	pCopyDstLayouts                                     &ImageLayout
	optimalTilingLayoutUUID                             [uuid_size]u8
	identicalMemoryTypeRequirements                     Bool32
}

// DeviceQueueGlobalPriorityCreateInfo extends VkDeviceQueueCreateInfo
pub type DeviceQueueGlobalPriorityCreateInfo = C.VkDeviceQueueGlobalPriorityCreateInfo

@[typedef]
pub struct C.VkDeviceQueueGlobalPriorityCreateInfo {
pub mut:
	sType          StructureType = StructureType.device_queue_global_priority_create_info
	pNext          voidptr       = unsafe { nil }
	globalPriority QueueGlobalPriority
}

// PhysicalDeviceGlobalPriorityQueryFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceGlobalPriorityQueryFeatures = C.VkPhysicalDeviceGlobalPriorityQueryFeatures

@[typedef]
pub struct C.VkPhysicalDeviceGlobalPriorityQueryFeatures {
pub mut:
	sType               StructureType = StructureType.physical_device_global_priority_query_features
	pNext               voidptr       = unsafe { nil }
	globalPriorityQuery Bool32
}

// QueueFamilyGlobalPriorityProperties extends VkQueueFamilyProperties2
pub type QueueFamilyGlobalPriorityProperties = C.VkQueueFamilyGlobalPriorityProperties

@[typedef]
pub struct C.VkQueueFamilyGlobalPriorityProperties {
pub mut:
	sType         StructureType = StructureType.queue_family_global_priority_properties
	pNext         voidptr       = unsafe { nil }
	priorityCount u32
	priorities    [max_global_priority_size]QueueGlobalPriority
}

// PhysicalDeviceIndexTypeUint8Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceIndexTypeUint8Features = C.VkPhysicalDeviceIndexTypeUint8Features

@[typedef]
pub struct C.VkPhysicalDeviceIndexTypeUint8Features {
pub mut:
	sType          StructureType = StructureType.physical_device_index_type_uint8_features
	pNext          voidptr       = unsafe { nil }
	indexTypeUint8 Bool32
}

pub type MemoryMapInfo = C.VkMemoryMapInfo

@[typedef]
pub struct C.VkMemoryMapInfo {
pub mut:
	sType  StructureType = StructureType.memory_map_info
	pNext  voidptr       = unsafe { nil }
	flags  MemoryMapFlags
	memory DeviceMemory
	offset DeviceSize
	size   DeviceSize
}

pub type MemoryUnmapInfo = C.VkMemoryUnmapInfo

@[typedef]
pub struct C.VkMemoryUnmapInfo {
pub mut:
	sType  StructureType = StructureType.memory_unmap_info
	pNext  voidptr       = unsafe { nil }
	flags  MemoryUnmapFlags
	memory DeviceMemory
}

// PhysicalDeviceMaintenance5Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMaintenance5Features = C.VkPhysicalDeviceMaintenance5Features

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance5Features {
pub mut:
	sType        StructureType = StructureType.physical_device_maintenance5_features
	pNext        voidptr       = unsafe { nil }
	maintenance5 Bool32
}

// PhysicalDeviceMaintenance5Properties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMaintenance5Properties = C.VkPhysicalDeviceMaintenance5Properties

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance5Properties {
pub mut:
	sType                                               StructureType = StructureType.physical_device_maintenance5_properties
	pNext                                               voidptr       = unsafe { nil }
	earlyFragmentMultisampleCoverageAfterSampleCounting Bool32
	earlyFragmentSampleMaskTestBeforeSampleCounting     Bool32
	depthStencilSwizzleOneSupport                       Bool32
	polygonModePointSize                                Bool32
	nonStrictSinglePixelWideLinesUseParallelogram       Bool32
	nonStrictWideLinesUseParallelogram                  Bool32
}

pub type ImageSubresource2 = C.VkImageSubresource2

@[typedef]
pub struct C.VkImageSubresource2 {
pub mut:
	sType            StructureType = StructureType.image_subresource2
	pNext            voidptr       = unsafe { nil }
	imageSubresource ImageSubresource
}

pub type DeviceImageSubresourceInfo = C.VkDeviceImageSubresourceInfo

@[typedef]
pub struct C.VkDeviceImageSubresourceInfo {
pub mut:
	sType        StructureType = StructureType.device_image_subresource_info
	pNext        voidptr       = unsafe { nil }
	pCreateInfo  &ImageCreateInfo
	pSubresource &ImageSubresource2
}

pub type SubresourceLayout2 = C.VkSubresourceLayout2

@[typedef]
pub struct C.VkSubresourceLayout2 {
pub mut:
	sType             StructureType = StructureType.subresource_layout2
	pNext             voidptr       = unsafe { nil }
	subresourceLayout SubresourceLayout
}

// BufferUsageFlags2CreateInfo extends VkBufferViewCreateInfo,VkBufferCreateInfo,VkPhysicalDeviceExternalBufferInfo,VkDescriptorBufferBindingInfoEXT
pub type BufferUsageFlags2CreateInfo = C.VkBufferUsageFlags2CreateInfo

@[typedef]
pub struct C.VkBufferUsageFlags2CreateInfo {
pub mut:
	sType StructureType = StructureType.buffer_usage_flags2_create_info
	pNext voidptr       = unsafe { nil }
	usage BufferUsageFlags2
}

// PhysicalDeviceMaintenance6Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMaintenance6Features = C.VkPhysicalDeviceMaintenance6Features

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance6Features {
pub mut:
	sType        StructureType = StructureType.physical_device_maintenance6_features
	pNext        voidptr       = unsafe { nil }
	maintenance6 Bool32
}

// PhysicalDeviceMaintenance6Properties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMaintenance6Properties = C.VkPhysicalDeviceMaintenance6Properties

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance6Properties {
pub mut:
	sType                                  StructureType = StructureType.physical_device_maintenance6_properties
	pNext                                  voidptr       = unsafe { nil }
	blockTexelViewCompatibleMultipleLayers Bool32
	maxCombinedImageSamplerDescriptorCount u32
	fragmentShadingRateClampCombinerInputs Bool32
}

// BindMemoryStatus extends VkBindBufferMemoryInfo,VkBindImageMemoryInfo
pub type BindMemoryStatus = C.VkBindMemoryStatus

@[typedef]
pub struct C.VkBindMemoryStatus {
pub mut:
	sType   StructureType = StructureType.bind_memory_status
	pNext   voidptr       = unsafe { nil }
	pResult &Result
}

// PhysicalDeviceHostImageCopyFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceHostImageCopyFeatures = C.VkPhysicalDeviceHostImageCopyFeatures

@[typedef]
pub struct C.VkPhysicalDeviceHostImageCopyFeatures {
pub mut:
	sType         StructureType = StructureType.physical_device_host_image_copy_features
	pNext         voidptr       = unsafe { nil }
	hostImageCopy Bool32
}

// PhysicalDeviceHostImageCopyProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceHostImageCopyProperties = C.VkPhysicalDeviceHostImageCopyProperties

@[typedef]
pub struct C.VkPhysicalDeviceHostImageCopyProperties {
pub mut:
	sType                           StructureType = StructureType.physical_device_host_image_copy_properties
	pNext                           voidptr       = unsafe { nil }
	copySrcLayoutCount              u32
	pCopySrcLayouts                 &ImageLayout
	copyDstLayoutCount              u32
	pCopyDstLayouts                 &ImageLayout
	optimalTilingLayoutUUID         [uuid_size]u8
	identicalMemoryTypeRequirements Bool32
}

pub type MemoryToImageCopy = C.VkMemoryToImageCopy

@[typedef]
pub struct C.VkMemoryToImageCopy {
pub mut:
	sType             StructureType = StructureType.memory_to_image_copy
	pNext             voidptr       = unsafe { nil }
	pHostPointer      voidptr
	memoryRowLength   u32
	memoryImageHeight u32
	imageSubresource  ImageSubresourceLayers
	imageOffset       Offset3D
	imageExtent       Extent3D
}

pub type ImageToMemoryCopy = C.VkImageToMemoryCopy

@[typedef]
pub struct C.VkImageToMemoryCopy {
pub mut:
	sType             StructureType = StructureType.image_to_memory_copy
	pNext             voidptr       = unsafe { nil }
	pHostPointer      voidptr
	memoryRowLength   u32
	memoryImageHeight u32
	imageSubresource  ImageSubresourceLayers
	imageOffset       Offset3D
	imageExtent       Extent3D
}

pub type CopyMemoryToImageInfo = C.VkCopyMemoryToImageInfo

@[typedef]
pub struct C.VkCopyMemoryToImageInfo {
pub mut:
	sType          StructureType = StructureType.copy_memory_to_image_info
	pNext          voidptr       = unsafe { nil }
	flags          HostImageCopyFlags
	dstImage       Image
	dstImageLayout ImageLayout
	regionCount    u32
	pRegions       &MemoryToImageCopy
}

pub type CopyImageToMemoryInfo = C.VkCopyImageToMemoryInfo

@[typedef]
pub struct C.VkCopyImageToMemoryInfo {
pub mut:
	sType          StructureType = StructureType.copy_image_to_memory_info
	pNext          voidptr       = unsafe { nil }
	flags          HostImageCopyFlags
	srcImage       Image
	srcImageLayout ImageLayout
	regionCount    u32
	pRegions       &ImageToMemoryCopy
}

pub type CopyImageToImageInfo = C.VkCopyImageToImageInfo

@[typedef]
pub struct C.VkCopyImageToImageInfo {
pub mut:
	sType          StructureType = StructureType.copy_image_to_image_info
	pNext          voidptr       = unsafe { nil }
	flags          HostImageCopyFlags
	srcImage       Image
	srcImageLayout ImageLayout
	dstImage       Image
	dstImageLayout ImageLayout
	regionCount    u32
	pRegions       &ImageCopy2
}

pub type HostImageLayoutTransitionInfo = C.VkHostImageLayoutTransitionInfo

@[typedef]
pub struct C.VkHostImageLayoutTransitionInfo {
pub mut:
	sType            StructureType = StructureType.host_image_layout_transition_info
	pNext            voidptr       = unsafe { nil }
	image            Image
	oldLayout        ImageLayout
	newLayout        ImageLayout
	subresourceRange ImageSubresourceRange
}

// SubresourceHostMemcpySize extends VkSubresourceLayout2
pub type SubresourceHostMemcpySize = C.VkSubresourceHostMemcpySize

@[typedef]
pub struct C.VkSubresourceHostMemcpySize {
pub mut:
	sType StructureType = StructureType.subresource_host_memcpy_size
	pNext voidptr       = unsafe { nil }
	size  DeviceSize
}

// HostImageCopyDevicePerformanceQuery extends VkImageFormatProperties2
pub type HostImageCopyDevicePerformanceQuery = C.VkHostImageCopyDevicePerformanceQuery

@[typedef]
pub struct C.VkHostImageCopyDevicePerformanceQuery {
pub mut:
	sType                 StructureType = StructureType.host_image_copy_device_performance_query
	pNext                 voidptr       = unsafe { nil }
	optimalDeviceAccess   Bool32
	identicalMemoryLayout Bool32
}

// PhysicalDeviceShaderSubgroupRotateFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderSubgroupRotateFeatures = C.VkPhysicalDeviceShaderSubgroupRotateFeatures

@[typedef]
pub struct C.VkPhysicalDeviceShaderSubgroupRotateFeatures {
pub mut:
	sType                         StructureType = StructureType.physical_device_shader_subgroup_rotate_features
	pNext                         voidptr       = unsafe { nil }
	shaderSubgroupRotate          Bool32
	shaderSubgroupRotateClustered Bool32
}

// PhysicalDeviceShaderFloatControls2Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderFloatControls2Features = C.VkPhysicalDeviceShaderFloatControls2Features

@[typedef]
pub struct C.VkPhysicalDeviceShaderFloatControls2Features {
pub mut:
	sType                StructureType = StructureType.physical_device_shader_float_controls2_features
	pNext                voidptr       = unsafe { nil }
	shaderFloatControls2 Bool32
}

// PhysicalDeviceShaderExpectAssumeFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderExpectAssumeFeatures = C.VkPhysicalDeviceShaderExpectAssumeFeatures

@[typedef]
pub struct C.VkPhysicalDeviceShaderExpectAssumeFeatures {
pub mut:
	sType              StructureType = StructureType.physical_device_shader_expect_assume_features
	pNext              voidptr       = unsafe { nil }
	shaderExpectAssume Bool32
}

// PipelineCreateFlags2CreateInfo extends VkComputePipelineCreateInfo,VkGraphicsPipelineCreateInfo,VkRayTracingPipelineCreateInfoNV,VkRayTracingPipelineCreateInfoKHR
pub type PipelineCreateFlags2CreateInfo = C.VkPipelineCreateFlags2CreateInfo

@[typedef]
pub struct C.VkPipelineCreateFlags2CreateInfo {
pub mut:
	sType StructureType = StructureType.pipeline_create_flags2_create_info
	pNext voidptr       = unsafe { nil }
	flags PipelineCreateFlags2
}

// PhysicalDevicePushDescriptorProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDevicePushDescriptorProperties = C.VkPhysicalDevicePushDescriptorProperties

@[typedef]
pub struct C.VkPhysicalDevicePushDescriptorProperties {
pub mut:
	sType              StructureType = StructureType.physical_device_push_descriptor_properties
	pNext              voidptr       = unsafe { nil }
	maxPushDescriptors u32
}

pub type BindDescriptorSetsInfo = C.VkBindDescriptorSetsInfo

@[typedef]
pub struct C.VkBindDescriptorSetsInfo {
pub mut:
	sType              StructureType = StructureType.bind_descriptor_sets_info
	pNext              voidptr       = unsafe { nil }
	stageFlags         ShaderStageFlags
	layout             PipelineLayout
	firstSet           u32
	descriptorSetCount u32
	pDescriptorSets    &DescriptorSet
	dynamicOffsetCount u32
	pDynamicOffsets    &u32
}

pub type PushConstantsInfo = C.VkPushConstantsInfo

@[typedef]
pub struct C.VkPushConstantsInfo {
pub mut:
	sType      StructureType = StructureType.push_constants_info
	pNext      voidptr       = unsafe { nil }
	layout     PipelineLayout
	stageFlags ShaderStageFlags
	offset     u32
	size       u32
	pValues    voidptr
}

pub type PushDescriptorSetInfo = C.VkPushDescriptorSetInfo

@[typedef]
pub struct C.VkPushDescriptorSetInfo {
pub mut:
	sType                StructureType = StructureType.push_descriptor_set_info
	pNext                voidptr       = unsafe { nil }
	stageFlags           ShaderStageFlags
	layout               PipelineLayout
	set                  u32
	descriptorWriteCount u32
	pDescriptorWrites    &WriteDescriptorSet
}

pub type PushDescriptorSetWithTemplateInfo = C.VkPushDescriptorSetWithTemplateInfo

@[typedef]
pub struct C.VkPushDescriptorSetWithTemplateInfo {
pub mut:
	sType                    StructureType = StructureType.push_descriptor_set_with_template_info
	pNext                    voidptr       = unsafe { nil }
	descriptorUpdateTemplate DescriptorUpdateTemplate
	layout                   PipelineLayout
	set                      u32
	pData                    voidptr
}

// PhysicalDevicePipelineProtectedAccessFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePipelineProtectedAccessFeatures = C.VkPhysicalDevicePipelineProtectedAccessFeatures

@[typedef]
pub struct C.VkPhysicalDevicePipelineProtectedAccessFeatures {
pub mut:
	sType                   StructureType = StructureType.physical_device_pipeline_protected_access_features
	pNext                   voidptr       = unsafe { nil }
	pipelineProtectedAccess Bool32
}

// PhysicalDevicePipelineRobustnessFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePipelineRobustnessFeatures = C.VkPhysicalDevicePipelineRobustnessFeatures

@[typedef]
pub struct C.VkPhysicalDevicePipelineRobustnessFeatures {
pub mut:
	sType              StructureType = StructureType.physical_device_pipeline_robustness_features
	pNext              voidptr       = unsafe { nil }
	pipelineRobustness Bool32
}

// PhysicalDevicePipelineRobustnessProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDevicePipelineRobustnessProperties = C.VkPhysicalDevicePipelineRobustnessProperties

@[typedef]
pub struct C.VkPhysicalDevicePipelineRobustnessProperties {
pub mut:
	sType                           StructureType = StructureType.physical_device_pipeline_robustness_properties
	pNext                           voidptr       = unsafe { nil }
	defaultRobustnessStorageBuffers PipelineRobustnessBufferBehavior
	defaultRobustnessUniformBuffers PipelineRobustnessBufferBehavior
	defaultRobustnessVertexInputs   PipelineRobustnessBufferBehavior
	defaultRobustnessImages         PipelineRobustnessImageBehavior
}

// PipelineRobustnessCreateInfo extends VkGraphicsPipelineCreateInfo,VkComputePipelineCreateInfo,VkPipelineShaderStageCreateInfo,VkRayTracingPipelineCreateInfoKHR
pub type PipelineRobustnessCreateInfo = C.VkPipelineRobustnessCreateInfo

@[typedef]
pub struct C.VkPipelineRobustnessCreateInfo {
pub mut:
	sType          StructureType = StructureType.pipeline_robustness_create_info
	pNext          voidptr       = unsafe { nil }
	storageBuffers PipelineRobustnessBufferBehavior
	uniformBuffers PipelineRobustnessBufferBehavior
	vertexInputs   PipelineRobustnessBufferBehavior
	images         PipelineRobustnessImageBehavior
}

// PhysicalDeviceLineRasterizationFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceLineRasterizationFeatures = C.VkPhysicalDeviceLineRasterizationFeatures

@[typedef]
pub struct C.VkPhysicalDeviceLineRasterizationFeatures {
pub mut:
	sType                    StructureType = StructureType.physical_device_line_rasterization_features
	pNext                    voidptr       = unsafe { nil }
	rectangularLines         Bool32
	bresenhamLines           Bool32
	smoothLines              Bool32
	stippledRectangularLines Bool32
	stippledBresenhamLines   Bool32
	stippledSmoothLines      Bool32
}

// PhysicalDeviceLineRasterizationProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceLineRasterizationProperties = C.VkPhysicalDeviceLineRasterizationProperties

@[typedef]
pub struct C.VkPhysicalDeviceLineRasterizationProperties {
pub mut:
	sType                     StructureType = StructureType.physical_device_line_rasterization_properties
	pNext                     voidptr       = unsafe { nil }
	lineSubPixelPrecisionBits u32
}

// PipelineRasterizationLineStateCreateInfo extends VkPipelineRasterizationStateCreateInfo
pub type PipelineRasterizationLineStateCreateInfo = C.VkPipelineRasterizationLineStateCreateInfo

@[typedef]
pub struct C.VkPipelineRasterizationLineStateCreateInfo {
pub mut:
	sType                 StructureType = StructureType.pipeline_rasterization_line_state_create_info
	pNext                 voidptr       = unsafe { nil }
	lineRasterizationMode LineRasterizationMode
	stippledLineEnable    Bool32
	lineStippleFactor     u32
	lineStipplePattern    u16
}

// PhysicalDeviceVertexAttributeDivisorProperties extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceVertexAttributeDivisorProperties = C.VkPhysicalDeviceVertexAttributeDivisorProperties

@[typedef]
pub struct C.VkPhysicalDeviceVertexAttributeDivisorProperties {
pub mut:
	sType                        StructureType = StructureType.physical_device_vertex_attribute_divisor_properties
	pNext                        voidptr       = unsafe { nil }
	maxVertexAttribDivisor       u32
	supportsNonZeroFirstInstance Bool32
}

pub type VertexInputBindingDivisorDescription = C.VkVertexInputBindingDivisorDescription

@[typedef]
pub struct C.VkVertexInputBindingDivisorDescription {
pub mut:
	binding u32
	divisor u32
}

// PipelineVertexInputDivisorStateCreateInfo extends VkPipelineVertexInputStateCreateInfo
pub type PipelineVertexInputDivisorStateCreateInfo = C.VkPipelineVertexInputDivisorStateCreateInfo

@[typedef]
pub struct C.VkPipelineVertexInputDivisorStateCreateInfo {
pub mut:
	sType                     StructureType = StructureType.pipeline_vertex_input_divisor_state_create_info
	pNext                     voidptr       = unsafe { nil }
	vertexBindingDivisorCount u32
	pVertexBindingDivisors    &VertexInputBindingDivisorDescription
}

// PhysicalDeviceVertexAttributeDivisorFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVertexAttributeDivisorFeatures = C.VkPhysicalDeviceVertexAttributeDivisorFeatures

@[typedef]
pub struct C.VkPhysicalDeviceVertexAttributeDivisorFeatures {
pub mut:
	sType                                  StructureType = StructureType.physical_device_vertex_attribute_divisor_features
	pNext                                  voidptr       = unsafe { nil }
	vertexAttributeInstanceRateDivisor     Bool32
	vertexAttributeInstanceRateZeroDivisor Bool32
}

pub type RenderingAreaInfo = C.VkRenderingAreaInfo

@[typedef]
pub struct C.VkRenderingAreaInfo {
pub mut:
	sType                   StructureType = StructureType.rendering_area_info
	pNext                   voidptr       = unsafe { nil }
	viewMask                u32
	colorAttachmentCount    u32
	pColorAttachmentFormats &Format
	depthAttachmentFormat   Format
	stencilAttachmentFormat Format
}

// PhysicalDeviceDynamicRenderingLocalReadFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDynamicRenderingLocalReadFeatures = C.VkPhysicalDeviceDynamicRenderingLocalReadFeatures

@[typedef]
pub struct C.VkPhysicalDeviceDynamicRenderingLocalReadFeatures {
pub mut:
	sType                     StructureType = StructureType.physical_device_dynamic_rendering_local_read_features
	pNext                     voidptr       = unsafe { nil }
	dynamicRenderingLocalRead Bool32
}

// RenderingAttachmentLocationInfo extends VkGraphicsPipelineCreateInfo,VkCommandBufferInheritanceInfo
pub type RenderingAttachmentLocationInfo = C.VkRenderingAttachmentLocationInfo

@[typedef]
pub struct C.VkRenderingAttachmentLocationInfo {
pub mut:
	sType                     StructureType = StructureType.rendering_attachment_location_info
	pNext                     voidptr       = unsafe { nil }
	colorAttachmentCount      u32
	pColorAttachmentLocations &u32
}

// RenderingInputAttachmentIndexInfo extends VkGraphicsPipelineCreateInfo,VkCommandBufferInheritanceInfo
pub type RenderingInputAttachmentIndexInfo = C.VkRenderingInputAttachmentIndexInfo

@[typedef]
pub struct C.VkRenderingInputAttachmentIndexInfo {
pub mut:
	sType                        StructureType = StructureType.rendering_input_attachment_index_info
	pNext                        voidptr       = unsafe { nil }
	colorAttachmentCount         u32
	pColorAttachmentInputIndices &u32
	pDepthInputAttachmentIndex   &u32
	pStencilInputAttachmentIndex &u32
}

@[keep_args_alive]
fn C.vkMapMemory2(device Device, p_memory_map_info &MemoryMapInfo, pp_data &voidptr) Result

pub type PFN_vkMapMemory2 = fn (device Device, p_memory_map_info &MemoryMapInfo, pp_data &voidptr) Result

@[inline]
pub fn map_memory2(device Device,
	p_memory_map_info &MemoryMapInfo,
	pp_data &voidptr) Result {
	return C.vkMapMemory2(device, p_memory_map_info, pp_data)
}

@[keep_args_alive]
fn C.vkUnmapMemory2(device Device, p_memory_unmap_info &MemoryUnmapInfo) Result

pub type PFN_vkUnmapMemory2 = fn (device Device, p_memory_unmap_info &MemoryUnmapInfo) Result

@[inline]
pub fn unmap_memory2(device Device,
	p_memory_unmap_info &MemoryUnmapInfo) Result {
	return C.vkUnmapMemory2(device, p_memory_unmap_info)
}

@[keep_args_alive]
fn C.vkGetDeviceImageSubresourceLayout(device Device, p_info &DeviceImageSubresourceInfo, mut p_layout SubresourceLayout2)

pub type PFN_vkGetDeviceImageSubresourceLayout = fn (device Device, p_info &DeviceImageSubresourceInfo, mut p_layout SubresourceLayout2)

@[inline]
pub fn get_device_image_subresource_layout(device Device,
	p_info &DeviceImageSubresourceInfo,
	mut p_layout SubresourceLayout2) {
	C.vkGetDeviceImageSubresourceLayout(device, p_info, mut p_layout)
}

@[keep_args_alive]
fn C.vkGetImageSubresourceLayout2(device Device, image Image, p_subresource &ImageSubresource2, mut p_layout SubresourceLayout2)

pub type PFN_vkGetImageSubresourceLayout2 = fn (device Device, image Image, p_subresource &ImageSubresource2, mut p_layout SubresourceLayout2)

@[inline]
pub fn get_image_subresource_layout2(device Device,
	image Image,
	p_subresource &ImageSubresource2,
	mut p_layout SubresourceLayout2) {
	C.vkGetImageSubresourceLayout2(device, image, p_subresource, mut p_layout)
}

@[keep_args_alive]
fn C.vkCopyMemoryToImage(device Device, p_copy_memory_to_image_info &CopyMemoryToImageInfo) Result

pub type PFN_vkCopyMemoryToImage = fn (device Device, p_copy_memory_to_image_info &CopyMemoryToImageInfo) Result

@[inline]
pub fn copy_memory_to_image(device Device,
	p_copy_memory_to_image_info &CopyMemoryToImageInfo) Result {
	return C.vkCopyMemoryToImage(device, p_copy_memory_to_image_info)
}

@[keep_args_alive]
fn C.vkCopyImageToMemory(device Device, p_copy_image_to_memory_info &CopyImageToMemoryInfo) Result

pub type PFN_vkCopyImageToMemory = fn (device Device, p_copy_image_to_memory_info &CopyImageToMemoryInfo) Result

@[inline]
pub fn copy_image_to_memory(device Device,
	p_copy_image_to_memory_info &CopyImageToMemoryInfo) Result {
	return C.vkCopyImageToMemory(device, p_copy_image_to_memory_info)
}

@[keep_args_alive]
fn C.vkCopyImageToImage(device Device, p_copy_image_to_image_info &CopyImageToImageInfo) Result

pub type PFN_vkCopyImageToImage = fn (device Device, p_copy_image_to_image_info &CopyImageToImageInfo) Result

@[inline]
pub fn copy_image_to_image(device Device,
	p_copy_image_to_image_info &CopyImageToImageInfo) Result {
	return C.vkCopyImageToImage(device, p_copy_image_to_image_info)
}

@[keep_args_alive]
fn C.vkTransitionImageLayout(device Device, transition_count u32, p_transitions &HostImageLayoutTransitionInfo) Result

pub type PFN_vkTransitionImageLayout = fn (device Device, transition_count u32, p_transitions &HostImageLayoutTransitionInfo) Result

@[inline]
pub fn transition_image_layout(device Device,
	transition_count u32,
	p_transitions &HostImageLayoutTransitionInfo) Result {
	return C.vkTransitionImageLayout(device, transition_count, p_transitions)
}

@[keep_args_alive]
fn C.vkCmdPushDescriptorSet(command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, layout PipelineLayout, set u32, descriptor_write_count u32, p_descriptor_writes &WriteDescriptorSet)

pub type PFN_vkCmdPushDescriptorSet = fn (command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, layout PipelineLayout, set u32, descriptor_write_count u32, p_descriptor_writes &WriteDescriptorSet)

@[inline]
pub fn cmd_push_descriptor_set(command_buffer CommandBuffer,
	pipeline_bind_point PipelineBindPoint,
	layout PipelineLayout,
	set u32,
	descriptor_write_count u32,
	p_descriptor_writes &WriteDescriptorSet) {
	C.vkCmdPushDescriptorSet(command_buffer, pipeline_bind_point, layout, set, descriptor_write_count,
		p_descriptor_writes)
}

@[keep_args_alive]
fn C.vkCmdPushDescriptorSetWithTemplate(command_buffer CommandBuffer, descriptor_update_template DescriptorUpdateTemplate, layout PipelineLayout, set u32, p_data voidptr)

pub type PFN_vkCmdPushDescriptorSetWithTemplate = fn (command_buffer CommandBuffer, descriptor_update_template DescriptorUpdateTemplate, layout PipelineLayout, set u32, p_data voidptr)

@[inline]
pub fn cmd_push_descriptor_set_with_template(command_buffer CommandBuffer,
	descriptor_update_template DescriptorUpdateTemplate,
	layout PipelineLayout,
	set u32,
	p_data voidptr) {
	C.vkCmdPushDescriptorSetWithTemplate(command_buffer, descriptor_update_template, layout,
		set, p_data)
}

@[keep_args_alive]
fn C.vkCmdBindDescriptorSets2(command_buffer CommandBuffer, p_bind_descriptor_sets_info &BindDescriptorSetsInfo)

pub type PFN_vkCmdBindDescriptorSets2 = fn (command_buffer CommandBuffer, p_bind_descriptor_sets_info &BindDescriptorSetsInfo)

@[inline]
pub fn cmd_bind_descriptor_sets2(command_buffer CommandBuffer,
	p_bind_descriptor_sets_info &BindDescriptorSetsInfo) {
	C.vkCmdBindDescriptorSets2(command_buffer, p_bind_descriptor_sets_info)
}

@[keep_args_alive]
fn C.vkCmdPushConstants2(command_buffer CommandBuffer, p_push_constants_info &PushConstantsInfo)

pub type PFN_vkCmdPushConstants2 = fn (command_buffer CommandBuffer, p_push_constants_info &PushConstantsInfo)

@[inline]
pub fn cmd_push_constants2(command_buffer CommandBuffer,
	p_push_constants_info &PushConstantsInfo) {
	C.vkCmdPushConstants2(command_buffer, p_push_constants_info)
}

@[keep_args_alive]
fn C.vkCmdPushDescriptorSet2(command_buffer CommandBuffer, p_push_descriptor_set_info &PushDescriptorSetInfo)

pub type PFN_vkCmdPushDescriptorSet2 = fn (command_buffer CommandBuffer, p_push_descriptor_set_info &PushDescriptorSetInfo)

@[inline]
pub fn cmd_push_descriptor_set2(command_buffer CommandBuffer,
	p_push_descriptor_set_info &PushDescriptorSetInfo) {
	C.vkCmdPushDescriptorSet2(command_buffer, p_push_descriptor_set_info)
}

@[keep_args_alive]
fn C.vkCmdPushDescriptorSetWithTemplate2(command_buffer CommandBuffer, p_push_descriptor_set_with_template_info &PushDescriptorSetWithTemplateInfo)

pub type PFN_vkCmdPushDescriptorSetWithTemplate2 = fn (command_buffer CommandBuffer, p_push_descriptor_set_with_template_info &PushDescriptorSetWithTemplateInfo)

@[inline]
pub fn cmd_push_descriptor_set_with_template2(command_buffer CommandBuffer,
	p_push_descriptor_set_with_template_info &PushDescriptorSetWithTemplateInfo) {
	C.vkCmdPushDescriptorSetWithTemplate2(command_buffer, p_push_descriptor_set_with_template_info)
}

@[keep_args_alive]
fn C.vkCmdSetLineStipple(command_buffer CommandBuffer, line_stipple_factor u32, line_stipple_pattern u16)

pub type PFN_vkCmdSetLineStipple = fn (command_buffer CommandBuffer, line_stipple_factor u32, line_stipple_pattern u16)

@[inline]
pub fn cmd_set_line_stipple(command_buffer CommandBuffer,
	line_stipple_factor u32,
	line_stipple_pattern u16) {
	C.vkCmdSetLineStipple(command_buffer, line_stipple_factor, line_stipple_pattern)
}

@[keep_args_alive]
fn C.vkCmdBindIndexBuffer2(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, size DeviceSize, index_type IndexType)

pub type PFN_vkCmdBindIndexBuffer2 = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, size DeviceSize, index_type IndexType)

@[inline]
pub fn cmd_bind_index_buffer2(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	size DeviceSize,
	index_type IndexType) {
	C.vkCmdBindIndexBuffer2(command_buffer, buffer, offset, size, index_type)
}

@[keep_args_alive]
fn C.vkGetRenderingAreaGranularity(device Device, p_rendering_area_info &RenderingAreaInfo, mut p_granularity Extent2D)

pub type PFN_vkGetRenderingAreaGranularity = fn (device Device, p_rendering_area_info &RenderingAreaInfo, mut p_granularity Extent2D)

@[inline]
pub fn get_rendering_area_granularity(device Device,
	p_rendering_area_info &RenderingAreaInfo,
	mut p_granularity Extent2D) {
	C.vkGetRenderingAreaGranularity(device, p_rendering_area_info, mut p_granularity)
}

@[keep_args_alive]
fn C.vkCmdSetRenderingAttachmentLocations(command_buffer CommandBuffer, p_location_info &RenderingAttachmentLocationInfo)

pub type PFN_vkCmdSetRenderingAttachmentLocations = fn (command_buffer CommandBuffer, p_location_info &RenderingAttachmentLocationInfo)

@[inline]
pub fn cmd_set_rendering_attachment_locations(command_buffer CommandBuffer,
	p_location_info &RenderingAttachmentLocationInfo) {
	C.vkCmdSetRenderingAttachmentLocations(command_buffer, p_location_info)
}

@[keep_args_alive]
fn C.vkCmdSetRenderingInputAttachmentIndices(command_buffer CommandBuffer, p_input_attachment_index_info &RenderingInputAttachmentIndexInfo)

pub type PFN_vkCmdSetRenderingInputAttachmentIndices = fn (command_buffer CommandBuffer, p_input_attachment_index_info &RenderingInputAttachmentIndexInfo)

@[inline]
pub fn cmd_set_rendering_input_attachment_indices(command_buffer CommandBuffer,
	p_input_attachment_index_info &RenderingInputAttachmentIndexInfo) {
	C.vkCmdSetRenderingInputAttachmentIndices(command_buffer, p_input_attachment_index_info)
}

// Pointer to VkSurfaceKHR_T
pub type SurfaceKHR = voidptr

pub const khr_surface_spec_version = 25
pub const khr_surface_extension_name = c'VK_KHR_surface'

pub enum PresentModeKHR as u32 {
	immediate                 = 0
	mailbox                   = 1
	fifo                      = 2
	fifo_relaxed              = 3
	shared_demand_refresh     = 1000111000
	shared_continuous_refresh = 1000111001
	fifo_latest_ready         = 1000361000
	max_enum_khr              = max_int
}

pub enum ColorSpaceKHR as u32 {
	srgb_nonlinear           = 0
	display_p3_nonlinear_ext = 1000104001
	extended_srgb_linear_ext = 1000104002
	display_p3_linear_ext    = 1000104003
	dci_p3_nonlinear_ext     = 1000104004
	bt709_linear_ext         = 1000104005
	bt709_nonlinear_ext      = 1000104006
	bt2020_linear_ext        = 1000104007
	hdr10_st2084_ext         = 1000104008
	// VK_COLOR_SPACE_DOLBYVISION_EXT is deprecated, but no reason was given in the API XML
	dolbyvision_ext             = 1000104009
	hdr10_hlg_ext               = 1000104010
	adobergb_linear_ext         = 1000104011
	adobergb_nonlinear_ext      = 1000104012
	pass_through_ext            = 1000104013
	extended_srgb_nonlinear_ext = 1000104014
	display_native_amd          = 1000213000
	max_enum_khr                = max_int
}

pub enum SurfaceTransformFlagBitsKHR as u32 {
	identity                    = u32(0x00000001)
	rotate90                    = u32(0x00000002)
	rotate180                   = u32(0x00000004)
	rotate270                   = u32(0x00000008)
	horizontal_mirror           = u32(0x00000010)
	horizontal_mirror_rotate90  = u32(0x00000020)
	horizontal_mirror_rotate180 = u32(0x00000040)
	horizontal_mirror_rotate270 = u32(0x00000080)
	inherit                     = u32(0x00000100)
	max_enum_khr                = max_int
}

pub enum CompositeAlphaFlagBitsKHR as u32 {
	opaque          = u32(0x00000001)
	pre_multiplied  = u32(0x00000002)
	post_multiplied = u32(0x00000004)
	inherit         = u32(0x00000008)
	max_enum_khr    = max_int
}
pub type CompositeAlphaFlagsKHR = u32
pub type SurfaceTransformFlagsKHR = u32
pub type SurfaceCapabilitiesKHR = C.VkSurfaceCapabilitiesKHR

@[typedef]
pub struct C.VkSurfaceCapabilitiesKHR {
pub mut:
	minImageCount           u32
	maxImageCount           u32
	currentExtent           Extent2D
	minImageExtent          Extent2D
	maxImageExtent          Extent2D
	maxImageArrayLayers     u32
	supportedTransforms     SurfaceTransformFlagsKHR
	currentTransform        SurfaceTransformFlagBitsKHR
	supportedCompositeAlpha CompositeAlphaFlagsKHR
	supportedUsageFlags     ImageUsageFlags
}

pub type SurfaceFormatKHR = C.VkSurfaceFormatKHR

@[typedef]
pub struct C.VkSurfaceFormatKHR {
pub mut:
	format     Format
	colorSpace ColorSpaceKHR
}

@[keep_args_alive]
fn C.vkDestroySurfaceKHR(instance Instance, surface SurfaceKHR, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroySurfaceKHR = fn (instance Instance, surface SurfaceKHR, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_surface_khr(instance Instance,
	surface SurfaceKHR,
	p_allocator &AllocationCallbacks) {
	C.vkDestroySurfaceKHR(instance, surface, p_allocator)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceSurfaceSupportKHR(physical_device PhysicalDevice, queue_family_index u32, surface SurfaceKHR, p_supported &Bool32) Result

pub type PFN_vkGetPhysicalDeviceSurfaceSupportKHR = fn (physical_device PhysicalDevice, queue_family_index u32, surface SurfaceKHR, p_supported &Bool32) Result

@[inline]
pub fn get_physical_device_surface_support_khr(physical_device PhysicalDevice,
	queue_family_index u32,
	surface SurfaceKHR,
	p_supported &Bool32) Result {
	return C.vkGetPhysicalDeviceSurfaceSupportKHR(physical_device, queue_family_index,
		surface, p_supported)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceSurfaceCapabilitiesKHR(physical_device PhysicalDevice, surface SurfaceKHR, mut p_surface_capabilities SurfaceCapabilitiesKHR) Result

pub type PFN_vkGetPhysicalDeviceSurfaceCapabilitiesKHR = fn (physical_device PhysicalDevice, surface SurfaceKHR, mut p_surface_capabilities SurfaceCapabilitiesKHR) Result

@[inline]
pub fn get_physical_device_surface_capabilities_khr(physical_device PhysicalDevice,
	surface SurfaceKHR,
	mut p_surface_capabilities SurfaceCapabilitiesKHR) Result {
	return C.vkGetPhysicalDeviceSurfaceCapabilitiesKHR(physical_device, surface, mut p_surface_capabilities)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceSurfaceFormatsKHR(physical_device PhysicalDevice, surface SurfaceKHR, p_surface_format_count &u32, mut p_surface_formats SurfaceFormatKHR) Result

pub type PFN_vkGetPhysicalDeviceSurfaceFormatsKHR = fn (physical_device PhysicalDevice, surface SurfaceKHR, p_surface_format_count &u32, mut p_surface_formats SurfaceFormatKHR) Result

@[inline]
pub fn get_physical_device_surface_formats_khr(physical_device PhysicalDevice,
	surface SurfaceKHR,
	p_surface_format_count &u32,
	mut p_surface_formats SurfaceFormatKHR) Result {
	return C.vkGetPhysicalDeviceSurfaceFormatsKHR(physical_device, surface, p_surface_format_count, mut
		p_surface_formats)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceSurfacePresentModesKHR(physical_device PhysicalDevice, surface SurfaceKHR, p_present_mode_count &u32, p_present_modes &PresentModeKHR) Result

pub type PFN_vkGetPhysicalDeviceSurfacePresentModesKHR = fn (physical_device PhysicalDevice, surface SurfaceKHR, p_present_mode_count &u32, p_present_modes &PresentModeKHR) Result

@[inline]
pub fn get_physical_device_surface_present_modes_khr(physical_device PhysicalDevice,
	surface SurfaceKHR,
	p_present_mode_count &u32,
	p_present_modes &PresentModeKHR) Result {
	return C.vkGetPhysicalDeviceSurfacePresentModesKHR(physical_device, surface, p_present_mode_count,
		p_present_modes)
}

// Pointer to VkSwapchainKHR_T
pub type SwapchainKHR = voidptr

pub const khr_swapchain_spec_version = 70
pub const khr_swapchain_extension_name = c'VK_KHR_swapchain'

pub enum SwapchainCreateFlagBitsKHR as u32 {
	split_instance_bind_regions = u32(0x00000001)
	protected                   = u32(0x00000002)
	mutable_format              = u32(0x00000004)
	present_id2                 = u32(0x00000040)
	present_wait2               = u32(0x00000080)
	deferred_memory_allocation  = u32(0x00000008)
	max_enum_khr                = max_int
}
pub type SwapchainCreateFlagsKHR = u32

pub enum DeviceGroupPresentModeFlagBitsKHR as u32 {
	local              = u32(0x00000001)
	remote             = u32(0x00000002)
	sum                = u32(0x00000004)
	local_multi_device = u32(0x00000008)
	max_enum_khr       = max_int
}
pub type DeviceGroupPresentModeFlagsKHR = u32
pub type SwapchainCreateInfoKHR = C.VkSwapchainCreateInfoKHR

@[typedef]
pub struct C.VkSwapchainCreateInfoKHR {
pub mut:
	sType                 StructureType = StructureType.swapchain_create_info_khr
	pNext                 voidptr       = unsafe { nil }
	flags                 SwapchainCreateFlagsKHR
	surface               SurfaceKHR
	minImageCount         u32
	imageFormat           Format
	imageColorSpace       ColorSpaceKHR
	imageExtent           Extent2D
	imageArrayLayers      u32
	imageUsage            ImageUsageFlags
	imageSharingMode      SharingMode
	queueFamilyIndexCount u32
	pQueueFamilyIndices   &u32
	preTransform          SurfaceTransformFlagBitsKHR
	compositeAlpha        CompositeAlphaFlagBitsKHR
	presentMode           PresentModeKHR
	clipped               Bool32
	oldSwapchain          SwapchainKHR
}

pub type PresentInfoKHR = C.VkPresentInfoKHR

@[typedef]
pub struct C.VkPresentInfoKHR {
pub mut:
	sType              StructureType = StructureType.present_info_khr
	pNext              voidptr       = unsafe { nil }
	waitSemaphoreCount u32
	pWaitSemaphores    &Semaphore
	swapchainCount     u32
	pSwapchains        &SwapchainKHR
	pImageIndices      &u32
	pResults           &Result
}

// ImageSwapchainCreateInfoKHR extends VkImageCreateInfo
pub type ImageSwapchainCreateInfoKHR = C.VkImageSwapchainCreateInfoKHR

@[typedef]
pub struct C.VkImageSwapchainCreateInfoKHR {
pub mut:
	sType     StructureType = StructureType.image_swapchain_create_info_khr
	pNext     voidptr       = unsafe { nil }
	swapchain SwapchainKHR
}

// BindImageMemorySwapchainInfoKHR extends VkBindImageMemoryInfo
pub type BindImageMemorySwapchainInfoKHR = C.VkBindImageMemorySwapchainInfoKHR

@[typedef]
pub struct C.VkBindImageMemorySwapchainInfoKHR {
pub mut:
	sType      StructureType = StructureType.bind_image_memory_swapchain_info_khr
	pNext      voidptr       = unsafe { nil }
	swapchain  SwapchainKHR
	imageIndex u32
}

pub type AcquireNextImageInfoKHR = C.VkAcquireNextImageInfoKHR

@[typedef]
pub struct C.VkAcquireNextImageInfoKHR {
pub mut:
	sType      StructureType = StructureType.acquire_next_image_info_khr
	pNext      voidptr       = unsafe { nil }
	swapchain  SwapchainKHR
	timeout    u64
	semaphore  Semaphore
	fence      Fence
	deviceMask u32
}

pub type DeviceGroupPresentCapabilitiesKHR = C.VkDeviceGroupPresentCapabilitiesKHR

@[typedef]
pub struct C.VkDeviceGroupPresentCapabilitiesKHR {
pub mut:
	sType       StructureType = StructureType.device_group_present_capabilities_khr
	pNext       voidptr       = unsafe { nil }
	presentMask [max_device_group_size]u32
	modes       DeviceGroupPresentModeFlagsKHR
}

// DeviceGroupPresentInfoKHR extends VkPresentInfoKHR
pub type DeviceGroupPresentInfoKHR = C.VkDeviceGroupPresentInfoKHR

@[typedef]
pub struct C.VkDeviceGroupPresentInfoKHR {
pub mut:
	sType          StructureType = StructureType.device_group_present_info_khr
	pNext          voidptr       = unsafe { nil }
	swapchainCount u32
	pDeviceMasks   &u32
	mode           DeviceGroupPresentModeFlagBitsKHR
}

// DeviceGroupSwapchainCreateInfoKHR extends VkSwapchainCreateInfoKHR
pub type DeviceGroupSwapchainCreateInfoKHR = C.VkDeviceGroupSwapchainCreateInfoKHR

@[typedef]
pub struct C.VkDeviceGroupSwapchainCreateInfoKHR {
pub mut:
	sType StructureType = StructureType.device_group_swapchain_create_info_khr
	pNext voidptr       = unsafe { nil }
	modes DeviceGroupPresentModeFlagsKHR
}

@[keep_args_alive]
fn C.vkCreateSwapchainKHR(device Device, p_create_info &SwapchainCreateInfoKHR, p_allocator &AllocationCallbacks, p_swapchain &SwapchainKHR) Result

pub type PFN_vkCreateSwapchainKHR = fn (device Device, p_create_info &SwapchainCreateInfoKHR, p_allocator &AllocationCallbacks, p_swapchain &SwapchainKHR) Result

@[inline]
pub fn create_swapchain_khr(device Device,
	p_create_info &SwapchainCreateInfoKHR,
	p_allocator &AllocationCallbacks,
	p_swapchain &SwapchainKHR) Result {
	return C.vkCreateSwapchainKHR(device, p_create_info, p_allocator, p_swapchain)
}

@[keep_args_alive]
fn C.vkDestroySwapchainKHR(device Device, swapchain SwapchainKHR, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroySwapchainKHR = fn (device Device, swapchain SwapchainKHR, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_swapchain_khr(device Device,
	swapchain SwapchainKHR,
	p_allocator &AllocationCallbacks) {
	C.vkDestroySwapchainKHR(device, swapchain, p_allocator)
}

@[keep_args_alive]
fn C.vkGetSwapchainImagesKHR(device Device, swapchain SwapchainKHR, p_swapchain_image_count &u32, p_swapchain_images &Image) Result

pub type PFN_vkGetSwapchainImagesKHR = fn (device Device, swapchain SwapchainKHR, p_swapchain_image_count &u32, p_swapchain_images &Image) Result

@[inline]
pub fn get_swapchain_images_khr(device Device,
	swapchain SwapchainKHR,
	p_swapchain_image_count &u32,
	p_swapchain_images &Image) Result {
	return C.vkGetSwapchainImagesKHR(device, swapchain, p_swapchain_image_count, p_swapchain_images)
}

@[keep_args_alive]
fn C.vkAcquireNextImageKHR(device Device, swapchain SwapchainKHR, timeout u64, semaphore Semaphore, fence Fence, p_image_index &u32) Result

pub type PFN_vkAcquireNextImageKHR = fn (device Device, swapchain SwapchainKHR, timeout u64, semaphore Semaphore, fence Fence, p_image_index &u32) Result

@[inline]
pub fn acquire_next_image_khr(device Device,
	swapchain SwapchainKHR,
	timeout u64,
	semaphore Semaphore,
	fence Fence,
	p_image_index &u32) Result {
	return C.vkAcquireNextImageKHR(device, swapchain, timeout, semaphore, fence, p_image_index)
}

@[keep_args_alive]
fn C.vkQueuePresentKHR(queue Queue, p_present_info &PresentInfoKHR) Result

pub type PFN_vkQueuePresentKHR = fn (queue Queue, p_present_info &PresentInfoKHR) Result

@[inline]
pub fn queue_present_khr(queue Queue,
	p_present_info &PresentInfoKHR) Result {
	return C.vkQueuePresentKHR(queue, p_present_info)
}

@[keep_args_alive]
fn C.vkGetDeviceGroupPresentCapabilitiesKHR(device Device, mut p_device_group_present_capabilities DeviceGroupPresentCapabilitiesKHR) Result

pub type PFN_vkGetDeviceGroupPresentCapabilitiesKHR = fn (device Device, mut p_device_group_present_capabilities DeviceGroupPresentCapabilitiesKHR) Result

@[inline]
pub fn get_device_group_present_capabilities_khr(device Device,
	mut p_device_group_present_capabilities DeviceGroupPresentCapabilitiesKHR) Result {
	return C.vkGetDeviceGroupPresentCapabilitiesKHR(device, mut p_device_group_present_capabilities)
}

@[keep_args_alive]
fn C.vkGetDeviceGroupSurfacePresentModesKHR(device Device, surface SurfaceKHR, p_modes &DeviceGroupPresentModeFlagsKHR) Result

pub type PFN_vkGetDeviceGroupSurfacePresentModesKHR = fn (device Device, surface SurfaceKHR, p_modes &DeviceGroupPresentModeFlagsKHR) Result

@[inline]
pub fn get_device_group_surface_present_modes_khr(device Device,
	surface SurfaceKHR,
	p_modes &DeviceGroupPresentModeFlagsKHR) Result {
	return C.vkGetDeviceGroupSurfacePresentModesKHR(device, surface, p_modes)
}

@[keep_args_alive]
fn C.vkGetPhysicalDevicePresentRectanglesKHR(physical_device PhysicalDevice, surface SurfaceKHR, p_rect_count &u32, mut p_rects Rect2D) Result

pub type PFN_vkGetPhysicalDevicePresentRectanglesKHR = fn (physical_device PhysicalDevice, surface SurfaceKHR, p_rect_count &u32, mut p_rects Rect2D) Result

@[inline]
pub fn get_physical_device_present_rectangles_khr(physical_device PhysicalDevice,
	surface SurfaceKHR,
	p_rect_count &u32,
	mut p_rects Rect2D) Result {
	return C.vkGetPhysicalDevicePresentRectanglesKHR(physical_device, surface, p_rect_count, mut
		p_rects)
}

@[keep_args_alive]
fn C.vkAcquireNextImage2KHR(device Device, p_acquire_info &AcquireNextImageInfoKHR, p_image_index &u32) Result

pub type PFN_vkAcquireNextImage2KHR = fn (device Device, p_acquire_info &AcquireNextImageInfoKHR, p_image_index &u32) Result

@[inline]
pub fn acquire_next_image2_khr(device Device,
	p_acquire_info &AcquireNextImageInfoKHR,
	p_image_index &u32) Result {
	return C.vkAcquireNextImage2KHR(device, p_acquire_info, p_image_index)
}

// Pointer to VkDisplayKHR_T
pub type DisplayKHR = voidptr

// Pointer to VkDisplayModeKHR_T
pub type DisplayModeKHR = voidptr

pub const khr_display_spec_version = 23
pub const khr_display_extension_name = c'VK_KHR_display'

pub type DisplayModeCreateFlagsKHR = u32

pub enum DisplayPlaneAlphaFlagBitsKHR as u32 {
	opaque                  = u32(0x00000001)
	global                  = u32(0x00000002)
	per_pixel               = u32(0x00000004)
	per_pixel_premultiplied = u32(0x00000008)
	max_enum_khr            = max_int
}
pub type DisplayPlaneAlphaFlagsKHR = u32
pub type DisplaySurfaceCreateFlagsKHR = u32
pub type DisplayModeParametersKHR = C.VkDisplayModeParametersKHR

@[typedef]
pub struct C.VkDisplayModeParametersKHR {
pub mut:
	visibleRegion Extent2D
	refreshRate   u32
}

pub type DisplayModeCreateInfoKHR = C.VkDisplayModeCreateInfoKHR

@[typedef]
pub struct C.VkDisplayModeCreateInfoKHR {
pub mut:
	sType      StructureType = StructureType.display_mode_create_info_khr
	pNext      voidptr       = unsafe { nil }
	flags      DisplayModeCreateFlagsKHR
	parameters DisplayModeParametersKHR
}

pub type DisplayModePropertiesKHR = C.VkDisplayModePropertiesKHR

@[typedef]
pub struct C.VkDisplayModePropertiesKHR {
pub mut:
	displayMode DisplayModeKHR
	parameters  DisplayModeParametersKHR
}

pub type DisplayPlaneCapabilitiesKHR = C.VkDisplayPlaneCapabilitiesKHR

@[typedef]
pub struct C.VkDisplayPlaneCapabilitiesKHR {
pub mut:
	supportedAlpha DisplayPlaneAlphaFlagsKHR
	minSrcPosition Offset2D
	maxSrcPosition Offset2D
	minSrcExtent   Extent2D
	maxSrcExtent   Extent2D
	minDstPosition Offset2D
	maxDstPosition Offset2D
	minDstExtent   Extent2D
	maxDstExtent   Extent2D
}

pub type DisplayPlanePropertiesKHR = C.VkDisplayPlanePropertiesKHR

@[typedef]
pub struct C.VkDisplayPlanePropertiesKHR {
pub mut:
	currentDisplay    DisplayKHR
	currentStackIndex u32
}

pub type DisplayPropertiesKHR = C.VkDisplayPropertiesKHR

@[typedef]
pub struct C.VkDisplayPropertiesKHR {
pub mut:
	display              DisplayKHR
	displayName          &char
	physicalDimensions   Extent2D
	physicalResolution   Extent2D
	supportedTransforms  SurfaceTransformFlagsKHR
	planeReorderPossible Bool32
	persistentContent    Bool32
}

pub type DisplaySurfaceCreateInfoKHR = C.VkDisplaySurfaceCreateInfoKHR

@[typedef]
pub struct C.VkDisplaySurfaceCreateInfoKHR {
pub mut:
	sType           StructureType = StructureType.display_surface_create_info_khr
	pNext           voidptr       = unsafe { nil }
	flags           DisplaySurfaceCreateFlagsKHR
	displayMode     DisplayModeKHR
	planeIndex      u32
	planeStackIndex u32
	transform       SurfaceTransformFlagBitsKHR
	globalAlpha     f32
	alphaMode       DisplayPlaneAlphaFlagBitsKHR
	imageExtent     Extent2D
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceDisplayPropertiesKHR(physical_device PhysicalDevice, p_property_count &u32, mut p_properties DisplayPropertiesKHR) Result

pub type PFN_vkGetPhysicalDeviceDisplayPropertiesKHR = fn (physical_device PhysicalDevice, p_property_count &u32, mut p_properties DisplayPropertiesKHR) Result

@[inline]
pub fn get_physical_device_display_properties_khr(physical_device PhysicalDevice,
	p_property_count &u32,
	mut p_properties DisplayPropertiesKHR) Result {
	return C.vkGetPhysicalDeviceDisplayPropertiesKHR(physical_device, p_property_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceDisplayPlanePropertiesKHR(physical_device PhysicalDevice, p_property_count &u32, mut p_properties DisplayPlanePropertiesKHR) Result

pub type PFN_vkGetPhysicalDeviceDisplayPlanePropertiesKHR = fn (physical_device PhysicalDevice, p_property_count &u32, mut p_properties DisplayPlanePropertiesKHR) Result

@[inline]
pub fn get_physical_device_display_plane_properties_khr(physical_device PhysicalDevice,
	p_property_count &u32,
	mut p_properties DisplayPlanePropertiesKHR) Result {
	return C.vkGetPhysicalDeviceDisplayPlanePropertiesKHR(physical_device, p_property_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkGetDisplayPlaneSupportedDisplaysKHR(physical_device PhysicalDevice, plane_index u32, p_display_count &u32, p_displays &DisplayKHR) Result

pub type PFN_vkGetDisplayPlaneSupportedDisplaysKHR = fn (physical_device PhysicalDevice, plane_index u32, p_display_count &u32, p_displays &DisplayKHR) Result

@[inline]
pub fn get_display_plane_supported_displays_khr(physical_device PhysicalDevice,
	plane_index u32,
	p_display_count &u32,
	p_displays &DisplayKHR) Result {
	return C.vkGetDisplayPlaneSupportedDisplaysKHR(physical_device, plane_index, p_display_count,
		p_displays)
}

@[keep_args_alive]
fn C.vkGetDisplayModePropertiesKHR(physical_device PhysicalDevice, display DisplayKHR, p_property_count &u32, mut p_properties DisplayModePropertiesKHR) Result

pub type PFN_vkGetDisplayModePropertiesKHR = fn (physical_device PhysicalDevice, display DisplayKHR, p_property_count &u32, mut p_properties DisplayModePropertiesKHR) Result

@[inline]
pub fn get_display_mode_properties_khr(physical_device PhysicalDevice,
	display DisplayKHR,
	p_property_count &u32,
	mut p_properties DisplayModePropertiesKHR) Result {
	return C.vkGetDisplayModePropertiesKHR(physical_device, display, p_property_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkCreateDisplayModeKHR(physical_device PhysicalDevice, display DisplayKHR, p_create_info &DisplayModeCreateInfoKHR, p_allocator &AllocationCallbacks, p_mode &DisplayModeKHR) Result

pub type PFN_vkCreateDisplayModeKHR = fn (physical_device PhysicalDevice, display DisplayKHR, p_create_info &DisplayModeCreateInfoKHR, p_allocator &AllocationCallbacks, p_mode &DisplayModeKHR) Result

@[inline]
pub fn create_display_mode_khr(physical_device PhysicalDevice,
	display DisplayKHR,
	p_create_info &DisplayModeCreateInfoKHR,
	p_allocator &AllocationCallbacks,
	p_mode &DisplayModeKHR) Result {
	return C.vkCreateDisplayModeKHR(physical_device, display, p_create_info, p_allocator,
		p_mode)
}

@[keep_args_alive]
fn C.vkGetDisplayPlaneCapabilitiesKHR(physical_device PhysicalDevice, mode DisplayModeKHR, plane_index u32, mut p_capabilities DisplayPlaneCapabilitiesKHR) Result

pub type PFN_vkGetDisplayPlaneCapabilitiesKHR = fn (physical_device PhysicalDevice, mode DisplayModeKHR, plane_index u32, mut p_capabilities DisplayPlaneCapabilitiesKHR) Result

@[inline]
pub fn get_display_plane_capabilities_khr(physical_device PhysicalDevice,
	mode DisplayModeKHR,
	plane_index u32,
	mut p_capabilities DisplayPlaneCapabilitiesKHR) Result {
	return C.vkGetDisplayPlaneCapabilitiesKHR(physical_device, mode, plane_index, mut
		p_capabilities)
}

@[keep_args_alive]
fn C.vkCreateDisplayPlaneSurfaceKHR(instance Instance, p_create_info &DisplaySurfaceCreateInfoKHR, p_allocator &AllocationCallbacks, p_surface &SurfaceKHR) Result

pub type PFN_vkCreateDisplayPlaneSurfaceKHR = fn (instance Instance, p_create_info &DisplaySurfaceCreateInfoKHR, p_allocator &AllocationCallbacks, p_surface &SurfaceKHR) Result

@[inline]
pub fn create_display_plane_surface_khr(instance Instance,
	p_create_info &DisplaySurfaceCreateInfoKHR,
	p_allocator &AllocationCallbacks,
	p_surface &SurfaceKHR) Result {
	return C.vkCreateDisplayPlaneSurfaceKHR(instance, p_create_info, p_allocator, p_surface)
}

pub const khr_display_swapchain_spec_version = 10
pub const khr_display_swapchain_extension_name = c'VK_KHR_display_swapchain'
// DisplayPresentInfoKHR extends VkPresentInfoKHR
pub type DisplayPresentInfoKHR = C.VkDisplayPresentInfoKHR

@[typedef]
pub struct C.VkDisplayPresentInfoKHR {
pub mut:
	sType      StructureType = StructureType.display_present_info_khr
	pNext      voidptr       = unsafe { nil }
	srcRect    Rect2D
	dstRect    Rect2D
	persistent Bool32
}

@[keep_args_alive]
fn C.vkCreateSharedSwapchainsKHR(device Device, swapchain_count u32, p_create_infos &SwapchainCreateInfoKHR, p_allocator &AllocationCallbacks, p_swapchains &SwapchainKHR) Result

pub type PFN_vkCreateSharedSwapchainsKHR = fn (device Device, swapchain_count u32, p_create_infos &SwapchainCreateInfoKHR, p_allocator &AllocationCallbacks, p_swapchains &SwapchainKHR) Result

@[inline]
pub fn create_shared_swapchains_khr(device Device,
	swapchain_count u32,
	p_create_infos &SwapchainCreateInfoKHR,
	p_allocator &AllocationCallbacks,
	p_swapchains &SwapchainKHR) Result {
	return C.vkCreateSharedSwapchainsKHR(device, swapchain_count, p_create_infos, p_allocator,
		p_swapchains)
}

pub const khr_sampler_mirror_clamp_to_edge_spec_version = 3
pub const khr_sampler_mirror_clamp_to_edge_extension_name = c'VK_KHR_sampler_mirror_clamp_to_edge'

// Pointer to VkVideoSessionKHR_T
pub type VideoSessionKHR = voidptr

// Pointer to VkVideoSessionParametersKHR_T
pub type VideoSessionParametersKHR = voidptr

pub const khr_video_queue_spec_version = 8
pub const khr_video_queue_extension_name = c'VK_KHR_video_queue'

pub enum QueryResultStatusKHR {
	error                               = -1
	not_ready                           = 0
	complete                            = 1
	insufficient_bitstream_buffer_range = -1000299000
	max_enum_khr                        = max_int
}

pub enum VideoCodecOperationFlagBitsKHR as u32 {
	none         = 0
	encode_h264  = u32(0x00010000)
	encode_h265  = u32(0x00020000)
	decode_h264  = u32(0x00000001)
	decode_h265  = u32(0x00000002)
	decode_av1   = u32(0x00000004)
	encode_av1   = u32(0x00040000)
	decode_vp9   = u32(0x00000008)
	max_enum_khr = max_int
}
pub type VideoCodecOperationFlagsKHR = u32

pub enum VideoChromaSubsamplingFlagBitsKHR as u32 {
	invalid      = 0
	monochrome   = u32(0x00000001)
	_420         = u32(0x00000002)
	_422         = u32(0x00000004)
	_444         = u32(0x00000008)
	max_enum_khr = max_int
}
pub type VideoChromaSubsamplingFlagsKHR = u32

pub enum VideoComponentBitDepthFlagBitsKHR as u32 {
	invalid      = 0
	_8           = u32(0x00000001)
	_10          = u32(0x00000004)
	_12          = u32(0x00000010)
	max_enum_khr = max_int
}
pub type VideoComponentBitDepthFlagsKHR = u32

pub enum VideoCapabilityFlagBitsKHR as u32 {
	protected_content         = u32(0x00000001)
	separate_reference_images = u32(0x00000002)
	max_enum_khr              = max_int
}
pub type VideoCapabilityFlagsKHR = u32

pub enum VideoSessionCreateFlagBitsKHR as u32 {
	protected_content                    = u32(0x00000001)
	allow_encode_parameter_optimizations = u32(0x00000002)
	inline_queries                       = u32(0x00000004)
	allow_encode_quantization_delta_map  = u32(0x00000008)
	allow_encode_emphasis_map            = u32(0x00000010)
	inline_session_parameters            = u32(0x00000020)
	max_enum_khr                         = max_int
}
pub type VideoSessionCreateFlagsKHR = u32

pub enum VideoSessionParametersCreateFlagBitsKHR as u32 {
	quantization_map_compatible = u32(0x00000001)
	max_enum_khr                = max_int
}
pub type VideoSessionParametersCreateFlagsKHR = u32
pub type VideoBeginCodingFlagsKHR = u32
pub type VideoEndCodingFlagsKHR = u32

pub enum VideoCodingControlFlagBitsKHR as u32 {
	reset                = u32(0x00000001)
	encode_rate_control  = u32(0x00000002)
	encode_quality_level = u32(0x00000004)
	max_enum_khr         = max_int
}
pub type VideoCodingControlFlagsKHR = u32

// QueueFamilyQueryResultStatusPropertiesKHR extends VkQueueFamilyProperties2
pub type QueueFamilyQueryResultStatusPropertiesKHR = C.VkQueueFamilyQueryResultStatusPropertiesKHR

@[typedef]
pub struct C.VkQueueFamilyQueryResultStatusPropertiesKHR {
pub mut:
	sType                    StructureType = StructureType.queue_family_query_result_status_properties_khr
	pNext                    voidptr       = unsafe { nil }
	queryResultStatusSupport Bool32
}

// QueueFamilyVideoPropertiesKHR extends VkQueueFamilyProperties2
pub type QueueFamilyVideoPropertiesKHR = C.VkQueueFamilyVideoPropertiesKHR

@[typedef]
pub struct C.VkQueueFamilyVideoPropertiesKHR {
pub mut:
	sType                StructureType = StructureType.queue_family_video_properties_khr
	pNext                voidptr       = unsafe { nil }
	videoCodecOperations VideoCodecOperationFlagsKHR
}

// VideoProfileInfoKHR extends VkQueryPoolCreateInfo
pub type VideoProfileInfoKHR = C.VkVideoProfileInfoKHR

@[typedef]
pub struct C.VkVideoProfileInfoKHR {
pub mut:
	sType               StructureType = StructureType.video_profile_info_khr
	pNext               voidptr       = unsafe { nil }
	videoCodecOperation VideoCodecOperationFlagBitsKHR
	chromaSubsampling   VideoChromaSubsamplingFlagsKHR
	lumaBitDepth        VideoComponentBitDepthFlagsKHR
	chromaBitDepth      VideoComponentBitDepthFlagsKHR
}

// VideoProfileListInfoKHR extends VkPhysicalDeviceImageFormatInfo2,VkPhysicalDeviceVideoFormatInfoKHR,VkImageCreateInfo,VkBufferCreateInfo
pub type VideoProfileListInfoKHR = C.VkVideoProfileListInfoKHR

@[typedef]
pub struct C.VkVideoProfileListInfoKHR {
pub mut:
	sType        StructureType = StructureType.video_profile_list_info_khr
	pNext        voidptr       = unsafe { nil }
	profileCount u32
	pProfiles    &VideoProfileInfoKHR
}

pub type VideoCapabilitiesKHR = C.VkVideoCapabilitiesKHR

@[typedef]
pub struct C.VkVideoCapabilitiesKHR {
pub mut:
	sType                             StructureType = StructureType.video_capabilities_khr
	pNext                             voidptr       = unsafe { nil }
	flags                             VideoCapabilityFlagsKHR
	minBitstreamBufferOffsetAlignment DeviceSize
	minBitstreamBufferSizeAlignment   DeviceSize
	pictureAccessGranularity          Extent2D
	minCodedExtent                    Extent2D
	maxCodedExtent                    Extent2D
	maxDpbSlots                       u32
	maxActiveReferencePictures        u32
	stdHeaderVersion                  ExtensionProperties
}

pub type PhysicalDeviceVideoFormatInfoKHR = C.VkPhysicalDeviceVideoFormatInfoKHR

@[typedef]
pub struct C.VkPhysicalDeviceVideoFormatInfoKHR {
pub mut:
	sType      StructureType = StructureType.physical_device_video_format_info_khr
	pNext      voidptr       = unsafe { nil }
	imageUsage ImageUsageFlags
}

pub type VideoFormatPropertiesKHR = C.VkVideoFormatPropertiesKHR

@[typedef]
pub struct C.VkVideoFormatPropertiesKHR {
pub mut:
	sType            StructureType = StructureType.video_format_properties_khr
	pNext            voidptr       = unsafe { nil }
	format           Format
	componentMapping ComponentMapping
	imageCreateFlags ImageCreateFlags
	imageType        ImageType
	imageTiling      ImageTiling
	imageUsageFlags  ImageUsageFlags
}

pub type VideoPictureResourceInfoKHR = C.VkVideoPictureResourceInfoKHR

@[typedef]
pub struct C.VkVideoPictureResourceInfoKHR {
pub mut:
	sType            StructureType = StructureType.video_picture_resource_info_khr
	pNext            voidptr       = unsafe { nil }
	codedOffset      Offset2D
	codedExtent      Extent2D
	baseArrayLayer   u32
	imageViewBinding ImageView
}

pub type VideoReferenceSlotInfoKHR = C.VkVideoReferenceSlotInfoKHR

@[typedef]
pub struct C.VkVideoReferenceSlotInfoKHR {
pub mut:
	sType            StructureType = StructureType.video_reference_slot_info_khr
	pNext            voidptr       = unsafe { nil }
	slotIndex        i32
	pPictureResource &VideoPictureResourceInfoKHR
}

pub type VideoSessionMemoryRequirementsKHR = C.VkVideoSessionMemoryRequirementsKHR

@[typedef]
pub struct C.VkVideoSessionMemoryRequirementsKHR {
pub mut:
	sType              StructureType = StructureType.video_session_memory_requirements_khr
	pNext              voidptr       = unsafe { nil }
	memoryBindIndex    u32
	memoryRequirements MemoryRequirements
}

pub type BindVideoSessionMemoryInfoKHR = C.VkBindVideoSessionMemoryInfoKHR

@[typedef]
pub struct C.VkBindVideoSessionMemoryInfoKHR {
pub mut:
	sType           StructureType = StructureType.bind_video_session_memory_info_khr
	pNext           voidptr       = unsafe { nil }
	memoryBindIndex u32
	memory          DeviceMemory
	memoryOffset    DeviceSize
	memorySize      DeviceSize
}

pub type VideoSessionCreateInfoKHR = C.VkVideoSessionCreateInfoKHR

@[typedef]
pub struct C.VkVideoSessionCreateInfoKHR {
pub mut:
	sType                      StructureType = StructureType.video_session_create_info_khr
	pNext                      voidptr       = unsafe { nil }
	queueFamilyIndex           u32
	flags                      VideoSessionCreateFlagsKHR
	pVideoProfile              &VideoProfileInfoKHR
	pictureFormat              Format
	maxCodedExtent             Extent2D
	referencePictureFormat     Format
	maxDpbSlots                u32
	maxActiveReferencePictures u32
	pStdHeaderVersion          &ExtensionProperties
}

pub type VideoSessionParametersCreateInfoKHR = C.VkVideoSessionParametersCreateInfoKHR

@[typedef]
pub struct C.VkVideoSessionParametersCreateInfoKHR {
pub mut:
	sType                          StructureType = StructureType.video_session_parameters_create_info_khr
	pNext                          voidptr       = unsafe { nil }
	flags                          VideoSessionParametersCreateFlagsKHR
	videoSessionParametersTemplate VideoSessionParametersKHR
	videoSession                   VideoSessionKHR
}

pub type VideoSessionParametersUpdateInfoKHR = C.VkVideoSessionParametersUpdateInfoKHR

@[typedef]
pub struct C.VkVideoSessionParametersUpdateInfoKHR {
pub mut:
	sType               StructureType = StructureType.video_session_parameters_update_info_khr
	pNext               voidptr       = unsafe { nil }
	updateSequenceCount u32
}

pub type VideoBeginCodingInfoKHR = C.VkVideoBeginCodingInfoKHR

@[typedef]
pub struct C.VkVideoBeginCodingInfoKHR {
pub mut:
	sType                  StructureType = StructureType.video_begin_coding_info_khr
	pNext                  voidptr       = unsafe { nil }
	flags                  VideoBeginCodingFlagsKHR
	videoSession           VideoSessionKHR
	videoSessionParameters VideoSessionParametersKHR
	referenceSlotCount     u32
	pReferenceSlots        &VideoReferenceSlotInfoKHR
}

pub type VideoEndCodingInfoKHR = C.VkVideoEndCodingInfoKHR

@[typedef]
pub struct C.VkVideoEndCodingInfoKHR {
pub mut:
	sType StructureType = StructureType.video_end_coding_info_khr
	pNext voidptr       = unsafe { nil }
	flags VideoEndCodingFlagsKHR
}

pub type VideoCodingControlInfoKHR = C.VkVideoCodingControlInfoKHR

@[typedef]
pub struct C.VkVideoCodingControlInfoKHR {
pub mut:
	sType StructureType = StructureType.video_coding_control_info_khr
	pNext voidptr       = unsafe { nil }
	flags VideoCodingControlFlagsKHR
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceVideoCapabilitiesKHR(physical_device PhysicalDevice, p_video_profile &VideoProfileInfoKHR, mut p_capabilities VideoCapabilitiesKHR) Result

pub type PFN_vkGetPhysicalDeviceVideoCapabilitiesKHR = fn (physical_device PhysicalDevice, p_video_profile &VideoProfileInfoKHR, mut p_capabilities VideoCapabilitiesKHR) Result

@[inline]
pub fn get_physical_device_video_capabilities_khr(physical_device PhysicalDevice,
	p_video_profile &VideoProfileInfoKHR,
	mut p_capabilities VideoCapabilitiesKHR) Result {
	return C.vkGetPhysicalDeviceVideoCapabilitiesKHR(physical_device, p_video_profile, mut
		p_capabilities)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceVideoFormatPropertiesKHR(physical_device PhysicalDevice, p_video_format_info &PhysicalDeviceVideoFormatInfoKHR, p_video_format_property_count &u32, mut p_video_format_properties VideoFormatPropertiesKHR) Result

pub type PFN_vkGetPhysicalDeviceVideoFormatPropertiesKHR = fn (physical_device PhysicalDevice, p_video_format_info &PhysicalDeviceVideoFormatInfoKHR, p_video_format_property_count &u32, mut p_video_format_properties VideoFormatPropertiesKHR) Result

@[inline]
pub fn get_physical_device_video_format_properties_khr(physical_device PhysicalDevice,
	p_video_format_info &PhysicalDeviceVideoFormatInfoKHR,
	p_video_format_property_count &u32,
	mut p_video_format_properties VideoFormatPropertiesKHR) Result {
	return C.vkGetPhysicalDeviceVideoFormatPropertiesKHR(physical_device, p_video_format_info,
		p_video_format_property_count, mut p_video_format_properties)
}

@[keep_args_alive]
fn C.vkCreateVideoSessionKHR(device Device, p_create_info &VideoSessionCreateInfoKHR, p_allocator &AllocationCallbacks, p_video_session &VideoSessionKHR) Result

pub type PFN_vkCreateVideoSessionKHR = fn (device Device, p_create_info &VideoSessionCreateInfoKHR, p_allocator &AllocationCallbacks, p_video_session &VideoSessionKHR) Result

@[inline]
pub fn create_video_session_khr(device Device,
	p_create_info &VideoSessionCreateInfoKHR,
	p_allocator &AllocationCallbacks,
	p_video_session &VideoSessionKHR) Result {
	return C.vkCreateVideoSessionKHR(device, p_create_info, p_allocator, p_video_session)
}

@[keep_args_alive]
fn C.vkDestroyVideoSessionKHR(device Device, video_session VideoSessionKHR, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyVideoSessionKHR = fn (device Device, video_session VideoSessionKHR, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_video_session_khr(device Device,
	video_session VideoSessionKHR,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyVideoSessionKHR(device, video_session, p_allocator)
}

@[keep_args_alive]
fn C.vkGetVideoSessionMemoryRequirementsKHR(device Device, video_session VideoSessionKHR, p_memory_requirements_count &u32, mut p_memory_requirements VideoSessionMemoryRequirementsKHR) Result

pub type PFN_vkGetVideoSessionMemoryRequirementsKHR = fn (device Device, video_session VideoSessionKHR, p_memory_requirements_count &u32, mut p_memory_requirements VideoSessionMemoryRequirementsKHR) Result

@[inline]
pub fn get_video_session_memory_requirements_khr(device Device,
	video_session VideoSessionKHR,
	p_memory_requirements_count &u32,
	mut p_memory_requirements VideoSessionMemoryRequirementsKHR) Result {
	return C.vkGetVideoSessionMemoryRequirementsKHR(device, video_session, p_memory_requirements_count, mut
		p_memory_requirements)
}

@[keep_args_alive]
fn C.vkBindVideoSessionMemoryKHR(device Device, video_session VideoSessionKHR, bind_session_memory_info_count u32, p_bind_session_memory_infos &BindVideoSessionMemoryInfoKHR) Result

pub type PFN_vkBindVideoSessionMemoryKHR = fn (device Device, video_session VideoSessionKHR, bind_session_memory_info_count u32, p_bind_session_memory_infos &BindVideoSessionMemoryInfoKHR) Result

@[inline]
pub fn bind_video_session_memory_khr(device Device,
	video_session VideoSessionKHR,
	bind_session_memory_info_count u32,
	p_bind_session_memory_infos &BindVideoSessionMemoryInfoKHR) Result {
	return C.vkBindVideoSessionMemoryKHR(device, video_session, bind_session_memory_info_count,
		p_bind_session_memory_infos)
}

@[keep_args_alive]
fn C.vkCreateVideoSessionParametersKHR(device Device, p_create_info &VideoSessionParametersCreateInfoKHR, p_allocator &AllocationCallbacks, p_video_session_parameters &VideoSessionParametersKHR) Result

pub type PFN_vkCreateVideoSessionParametersKHR = fn (device Device, p_create_info &VideoSessionParametersCreateInfoKHR, p_allocator &AllocationCallbacks, p_video_session_parameters &VideoSessionParametersKHR) Result

@[inline]
pub fn create_video_session_parameters_khr(device Device,
	p_create_info &VideoSessionParametersCreateInfoKHR,
	p_allocator &AllocationCallbacks,
	p_video_session_parameters &VideoSessionParametersKHR) Result {
	return C.vkCreateVideoSessionParametersKHR(device, p_create_info, p_allocator, p_video_session_parameters)
}

@[keep_args_alive]
fn C.vkUpdateVideoSessionParametersKHR(device Device, video_session_parameters VideoSessionParametersKHR, p_update_info &VideoSessionParametersUpdateInfoKHR) Result

pub type PFN_vkUpdateVideoSessionParametersKHR = fn (device Device, video_session_parameters VideoSessionParametersKHR, p_update_info &VideoSessionParametersUpdateInfoKHR) Result

@[inline]
pub fn update_video_session_parameters_khr(device Device,
	video_session_parameters VideoSessionParametersKHR,
	p_update_info &VideoSessionParametersUpdateInfoKHR) Result {
	return C.vkUpdateVideoSessionParametersKHR(device, video_session_parameters, p_update_info)
}

@[keep_args_alive]
fn C.vkDestroyVideoSessionParametersKHR(device Device, video_session_parameters VideoSessionParametersKHR, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyVideoSessionParametersKHR = fn (device Device, video_session_parameters VideoSessionParametersKHR, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_video_session_parameters_khr(device Device,
	video_session_parameters VideoSessionParametersKHR,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyVideoSessionParametersKHR(device, video_session_parameters, p_allocator)
}

@[keep_args_alive]
fn C.vkCmdBeginVideoCodingKHR(command_buffer CommandBuffer, p_begin_info &VideoBeginCodingInfoKHR)

pub type PFN_vkCmdBeginVideoCodingKHR = fn (command_buffer CommandBuffer, p_begin_info &VideoBeginCodingInfoKHR)

@[inline]
pub fn cmd_begin_video_coding_khr(command_buffer CommandBuffer,
	p_begin_info &VideoBeginCodingInfoKHR) {
	C.vkCmdBeginVideoCodingKHR(command_buffer, p_begin_info)
}

@[keep_args_alive]
fn C.vkCmdEndVideoCodingKHR(command_buffer CommandBuffer, p_end_coding_info &VideoEndCodingInfoKHR)

pub type PFN_vkCmdEndVideoCodingKHR = fn (command_buffer CommandBuffer, p_end_coding_info &VideoEndCodingInfoKHR)

@[inline]
pub fn cmd_end_video_coding_khr(command_buffer CommandBuffer,
	p_end_coding_info &VideoEndCodingInfoKHR) {
	C.vkCmdEndVideoCodingKHR(command_buffer, p_end_coding_info)
}

@[keep_args_alive]
fn C.vkCmdControlVideoCodingKHR(command_buffer CommandBuffer, p_coding_control_info &VideoCodingControlInfoKHR)

pub type PFN_vkCmdControlVideoCodingKHR = fn (command_buffer CommandBuffer, p_coding_control_info &VideoCodingControlInfoKHR)

@[inline]
pub fn cmd_control_video_coding_khr(command_buffer CommandBuffer,
	p_coding_control_info &VideoCodingControlInfoKHR) {
	C.vkCmdControlVideoCodingKHR(command_buffer, p_coding_control_info)
}

pub const khr_video_decode_queue_spec_version = 8
pub const khr_video_decode_queue_extension_name = c'VK_KHR_video_decode_queue'

pub enum VideoDecodeCapabilityFlagBitsKHR as u32 {
	dpb_and_output_coincide = u32(0x00000001)
	dpb_and_output_distinct = u32(0x00000002)
	max_enum_khr            = max_int
}
pub type VideoDecodeCapabilityFlagsKHR = u32

pub enum VideoDecodeUsageFlagBitsKHR as u32 {
	default      = 0
	transcoding  = u32(0x00000001)
	offline      = u32(0x00000002)
	streaming    = u32(0x00000004)
	max_enum_khr = max_int
}
pub type VideoDecodeUsageFlagsKHR = u32
pub type VideoDecodeFlagsKHR = u32

// VideoDecodeCapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoDecodeCapabilitiesKHR = C.VkVideoDecodeCapabilitiesKHR

@[typedef]
pub struct C.VkVideoDecodeCapabilitiesKHR {
pub mut:
	sType StructureType = StructureType.video_decode_capabilities_khr
	pNext voidptr       = unsafe { nil }
	flags VideoDecodeCapabilityFlagsKHR
}

// VideoDecodeUsageInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub type VideoDecodeUsageInfoKHR = C.VkVideoDecodeUsageInfoKHR

@[typedef]
pub struct C.VkVideoDecodeUsageInfoKHR {
pub mut:
	sType           StructureType = StructureType.video_decode_usage_info_khr
	pNext           voidptr       = unsafe { nil }
	videoUsageHints VideoDecodeUsageFlagsKHR
}

pub type VideoDecodeInfoKHR = C.VkVideoDecodeInfoKHR

@[typedef]
pub struct C.VkVideoDecodeInfoKHR {
pub mut:
	sType               StructureType = StructureType.video_decode_info_khr
	pNext               voidptr       = unsafe { nil }
	flags               VideoDecodeFlagsKHR
	srcBuffer           Buffer
	srcBufferOffset     DeviceSize
	srcBufferRange      DeviceSize
	dstPictureResource  VideoPictureResourceInfoKHR
	pSetupReferenceSlot &VideoReferenceSlotInfoKHR
	referenceSlotCount  u32
	pReferenceSlots     &VideoReferenceSlotInfoKHR
}

@[keep_args_alive]
fn C.vkCmdDecodeVideoKHR(command_buffer CommandBuffer, p_decode_info &VideoDecodeInfoKHR)

pub type PFN_vkCmdDecodeVideoKHR = fn (command_buffer CommandBuffer, p_decode_info &VideoDecodeInfoKHR)

@[inline]
pub fn cmd_decode_video_khr(command_buffer CommandBuffer,
	p_decode_info &VideoDecodeInfoKHR) {
	C.vkCmdDecodeVideoKHR(command_buffer, p_decode_info)
}

pub const khr_video_encode_h264_spec_version = 14
pub const khr_video_encode_h264_extension_name = c'VK_KHR_video_encode_h264'

pub enum VideoEncodeH264CapabilityFlagBitsKHR as u32 {
	hrd_compliance                    = u32(0x00000001)
	prediction_weight_table_generated = u32(0x00000002)
	row_unaligned_slice               = u32(0x00000004)
	different_slice_type              = u32(0x00000008)
	b_frame_in_l0_list                = u32(0x00000010)
	b_frame_in_l1_list                = u32(0x00000020)
	per_picture_type_min_max_qp       = u32(0x00000040)
	per_slice_constant_qp             = u32(0x00000080)
	generate_prefix_nalu              = u32(0x00000100)
	b_picture_intra_refresh           = u32(0x00000400)
	mb_qp_diff_wraparound             = u32(0x00000200)
	max_enum_khr                      = max_int
}
pub type VideoEncodeH264CapabilityFlagsKHR = u32

pub enum VideoEncodeH264StdFlagBitsKHR as u32 {
	separate_color_plane_flag_set            = u32(0x00000001)
	qpprime_y_zero_transform_bypass_flag_set = u32(0x00000002)
	scaling_matrix_present_flag_set          = u32(0x00000004)
	chroma_qp_index_offset                   = u32(0x00000008)
	second_chroma_qp_index_offset            = u32(0x00000010)
	pic_init_qp_minus26                      = u32(0x00000020)
	weighted_pred_flag_set                   = u32(0x00000040)
	weighted_bipred_idc_explicit             = u32(0x00000080)
	weighted_bipred_idc_implicit             = u32(0x00000100)
	transform8x8_mode_flag_set               = u32(0x00000200)
	direct_spatial_mv_pred_flag_unset        = u32(0x00000400)
	entropy_coding_mode_flag_unset           = u32(0x00000800)
	entropy_coding_mode_flag_set             = u32(0x00001000)
	direct8x8_inference_flag_unset           = u32(0x00002000)
	constrained_intra_pred_flag_set          = u32(0x00004000)
	deblocking_filter_disabled               = u32(0x00008000)
	deblocking_filter_enabled                = u32(0x00010000)
	deblocking_filter_partial                = u32(0x00020000)
	slice_qp_delta                           = u32(0x00080000)
	different_slice_qp_delta                 = u32(0x00100000)
	max_enum_khr                             = max_int
}
pub type VideoEncodeH264StdFlagsKHR = u32

pub enum VideoEncodeH264RateControlFlagBitsKHR as u32 {
	attempt_hrd_compliance        = u32(0x00000001)
	regular_gop                   = u32(0x00000002)
	reference_pattern_flat        = u32(0x00000004)
	reference_pattern_dyadic      = u32(0x00000008)
	temporal_layer_pattern_dyadic = u32(0x00000010)
	max_enum_khr                  = max_int
}
pub type VideoEncodeH264RateControlFlagsKHR = u32

// VideoEncodeH264CapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoEncodeH264CapabilitiesKHR = C.VkVideoEncodeH264CapabilitiesKHR

@[typedef]
pub struct C.VkVideoEncodeH264CapabilitiesKHR {
pub mut:
	sType                            StructureType = StructureType.video_encode_h264_capabilities_khr
	pNext                            voidptr       = unsafe { nil }
	flags                            VideoEncodeH264CapabilityFlagsKHR
	maxLevelIdc                      StdVideoH264LevelIdc
	maxSliceCount                    u32
	maxPPictureL0ReferenceCount      u32
	maxBPictureL0ReferenceCount      u32
	maxL1ReferenceCount              u32
	maxTemporalLayerCount            u32
	expectDyadicTemporalLayerPattern Bool32
	minQp                            i32
	maxQp                            i32
	prefersGopRemainingFrames        Bool32
	requiresGopRemainingFrames       Bool32
	stdSyntaxFlags                   VideoEncodeH264StdFlagsKHR
}

pub type VideoEncodeH264QpKHR = C.VkVideoEncodeH264QpKHR

@[typedef]
pub struct C.VkVideoEncodeH264QpKHR {
pub mut:
	qpI i32
	qpP i32
	qpB i32
}

// VideoEncodeH264QualityLevelPropertiesKHR extends VkVideoEncodeQualityLevelPropertiesKHR
pub type VideoEncodeH264QualityLevelPropertiesKHR = C.VkVideoEncodeH264QualityLevelPropertiesKHR

@[typedef]
pub struct C.VkVideoEncodeH264QualityLevelPropertiesKHR {
pub mut:
	sType                             StructureType = StructureType.video_encode_h264_quality_level_properties_khr
	pNext                             voidptr       = unsafe { nil }
	preferredRateControlFlags         VideoEncodeH264RateControlFlagsKHR
	preferredGopFrameCount            u32
	preferredIdrPeriod                u32
	preferredConsecutiveBFrameCount   u32
	preferredTemporalLayerCount       u32
	preferredConstantQp               VideoEncodeH264QpKHR
	preferredMaxL0ReferenceCount      u32
	preferredMaxL1ReferenceCount      u32
	preferredStdEntropyCodingModeFlag Bool32
}

// VideoEncodeH264SessionCreateInfoKHR extends VkVideoSessionCreateInfoKHR
pub type VideoEncodeH264SessionCreateInfoKHR = C.VkVideoEncodeH264SessionCreateInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264SessionCreateInfoKHR {
pub mut:
	sType          StructureType = StructureType.video_encode_h264_session_create_info_khr
	pNext          voidptr       = unsafe { nil }
	useMaxLevelIdc Bool32
	maxLevelIdc    StdVideoH264LevelIdc
}

// VideoEncodeH264SessionParametersAddInfoKHR extends VkVideoSessionParametersUpdateInfoKHR
pub type VideoEncodeH264SessionParametersAddInfoKHR = C.VkVideoEncodeH264SessionParametersAddInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264SessionParametersAddInfoKHR {
pub mut:
	sType       StructureType = StructureType.video_encode_h264_session_parameters_add_info_khr
	pNext       voidptr       = unsafe { nil }
	stdSPSCount u32
	pStdSPSs    &StdVideoH264SequenceParameterSet
	stdPPSCount u32
	pStdPPSs    &StdVideoH264PictureParameterSet
}

// VideoEncodeH264SessionParametersCreateInfoKHR extends VkVideoSessionParametersCreateInfoKHR
pub type VideoEncodeH264SessionParametersCreateInfoKHR = C.VkVideoEncodeH264SessionParametersCreateInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264SessionParametersCreateInfoKHR {
pub mut:
	sType              StructureType = StructureType.video_encode_h264_session_parameters_create_info_khr
	pNext              voidptr       = unsafe { nil }
	maxStdSPSCount     u32
	maxStdPPSCount     u32
	pParametersAddInfo &VideoEncodeH264SessionParametersAddInfoKHR
}

// VideoEncodeH264SessionParametersGetInfoKHR extends VkVideoEncodeSessionParametersGetInfoKHR
pub type VideoEncodeH264SessionParametersGetInfoKHR = C.VkVideoEncodeH264SessionParametersGetInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264SessionParametersGetInfoKHR {
pub mut:
	sType       StructureType = StructureType.video_encode_h264_session_parameters_get_info_khr
	pNext       voidptr       = unsafe { nil }
	writeStdSPS Bool32
	writeStdPPS Bool32
	stdSPSId    u32
	stdPPSId    u32
}

// VideoEncodeH264SessionParametersFeedbackInfoKHR extends VkVideoEncodeSessionParametersFeedbackInfoKHR
pub type VideoEncodeH264SessionParametersFeedbackInfoKHR = C.VkVideoEncodeH264SessionParametersFeedbackInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264SessionParametersFeedbackInfoKHR {
pub mut:
	sType              StructureType = StructureType.video_encode_h264_session_parameters_feedback_info_khr
	pNext              voidptr       = unsafe { nil }
	hasStdSPSOverrides Bool32
	hasStdPPSOverrides Bool32
}

pub type VideoEncodeH264NaluSliceInfoKHR = C.VkVideoEncodeH264NaluSliceInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264NaluSliceInfoKHR {
pub mut:
	sType           StructureType = StructureType.video_encode_h264_nalu_slice_info_khr
	pNext           voidptr       = unsafe { nil }
	constantQp      i32
	pStdSliceHeader &StdVideoEncodeH264SliceHeader
}

// VideoEncodeH264PictureInfoKHR extends VkVideoEncodeInfoKHR
pub type VideoEncodeH264PictureInfoKHR = C.VkVideoEncodeH264PictureInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264PictureInfoKHR {
pub mut:
	sType               StructureType = StructureType.video_encode_h264_picture_info_khr
	pNext               voidptr       = unsafe { nil }
	naluSliceEntryCount u32
	pNaluSliceEntries   &VideoEncodeH264NaluSliceInfoKHR
	pStdPictureInfo     &StdVideoEncodeH264PictureInfo
	generatePrefixNalu  Bool32
}

// VideoEncodeH264DpbSlotInfoKHR extends VkVideoReferenceSlotInfoKHR
pub type VideoEncodeH264DpbSlotInfoKHR = C.VkVideoEncodeH264DpbSlotInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264DpbSlotInfoKHR {
pub mut:
	sType             StructureType = StructureType.video_encode_h264_dpb_slot_info_khr
	pNext             voidptr       = unsafe { nil }
	pStdReferenceInfo &StdVideoEncodeH264ReferenceInfo
}

// VideoEncodeH264ProfileInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub type VideoEncodeH264ProfileInfoKHR = C.VkVideoEncodeH264ProfileInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264ProfileInfoKHR {
pub mut:
	sType         StructureType = StructureType.video_encode_h264_profile_info_khr
	pNext         voidptr       = unsafe { nil }
	stdProfileIdc StdVideoH264ProfileIdc
}

// VideoEncodeH264RateControlInfoKHR extends VkVideoCodingControlInfoKHR,VkVideoBeginCodingInfoKHR
pub type VideoEncodeH264RateControlInfoKHR = C.VkVideoEncodeH264RateControlInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264RateControlInfoKHR {
pub mut:
	sType                  StructureType = StructureType.video_encode_h264_rate_control_info_khr
	pNext                  voidptr       = unsafe { nil }
	flags                  VideoEncodeH264RateControlFlagsKHR
	gopFrameCount          u32
	idrPeriod              u32
	consecutiveBFrameCount u32
	temporalLayerCount     u32
}

pub type VideoEncodeH264FrameSizeKHR = C.VkVideoEncodeH264FrameSizeKHR

@[typedef]
pub struct C.VkVideoEncodeH264FrameSizeKHR {
pub mut:
	frameISize u32
	framePSize u32
	frameBSize u32
}

// VideoEncodeH264RateControlLayerInfoKHR extends VkVideoEncodeRateControlLayerInfoKHR
pub type VideoEncodeH264RateControlLayerInfoKHR = C.VkVideoEncodeH264RateControlLayerInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264RateControlLayerInfoKHR {
pub mut:
	sType           StructureType = StructureType.video_encode_h264_rate_control_layer_info_khr
	pNext           voidptr       = unsafe { nil }
	useMinQp        Bool32
	minQp           VideoEncodeH264QpKHR
	useMaxQp        Bool32
	maxQp           VideoEncodeH264QpKHR
	useMaxFrameSize Bool32
	maxFrameSize    VideoEncodeH264FrameSizeKHR
}

// VideoEncodeH264GopRemainingFrameInfoKHR extends VkVideoBeginCodingInfoKHR
pub type VideoEncodeH264GopRemainingFrameInfoKHR = C.VkVideoEncodeH264GopRemainingFrameInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH264GopRemainingFrameInfoKHR {
pub mut:
	sType                 StructureType = StructureType.video_encode_h264_gop_remaining_frame_info_khr
	pNext                 voidptr       = unsafe { nil }
	useGopRemainingFrames Bool32
	gopRemainingI         u32
	gopRemainingP         u32
	gopRemainingB         u32
}

pub const khr_video_encode_h265_spec_version = 14
pub const khr_video_encode_h265_extension_name = c'VK_KHR_video_encode_h265'

pub enum VideoEncodeH265CapabilityFlagBitsKHR as u32 {
	hrd_compliance                    = u32(0x00000001)
	prediction_weight_table_generated = u32(0x00000002)
	row_unaligned_slice_segment       = u32(0x00000004)
	different_slice_segment_type      = u32(0x00000008)
	b_frame_in_l0_list                = u32(0x00000010)
	b_frame_in_l1_list                = u32(0x00000020)
	per_picture_type_min_max_qp       = u32(0x00000040)
	per_slice_segment_constant_qp     = u32(0x00000080)
	multiple_tiles_per_slice_segment  = u32(0x00000100)
	multiple_slice_segments_per_tile  = u32(0x00000200)
	b_picture_intra_refresh           = u32(0x00000800)
	cu_qp_diff_wraparound             = u32(0x00000400)
	max_enum_khr                      = max_int
}
pub type VideoEncodeH265CapabilityFlagsKHR = u32

pub enum VideoEncodeH265StdFlagBitsKHR as u32 {
	separate_color_plane_flag_set                = u32(0x00000001)
	sample_adaptive_offset_enabled_flag_set      = u32(0x00000002)
	scaling_list_data_present_flag_set           = u32(0x00000004)
	pcm_enabled_flag_set                         = u32(0x00000008)
	sps_temporal_mvp_enabled_flag_set            = u32(0x00000010)
	init_qp_minus26                              = u32(0x00000020)
	weighted_pred_flag_set                       = u32(0x00000040)
	weighted_bipred_flag_set                     = u32(0x00000080)
	log2_parallel_merge_level_minus2             = u32(0x00000100)
	sign_data_hiding_enabled_flag_set            = u32(0x00000200)
	transform_skip_enabled_flag_set              = u32(0x00000400)
	transform_skip_enabled_flag_unset            = u32(0x00000800)
	pps_slice_chroma_qp_offsets_present_flag_set = u32(0x00001000)
	transquant_bypass_enabled_flag_set           = u32(0x00002000)
	constrained_intra_pred_flag_set              = u32(0x00004000)
	entropy_coding_sync_enabled_flag_set         = u32(0x00008000)
	deblocking_filter_override_enabled_flag_set  = u32(0x00010000)
	dependent_slice_segments_enabled_flag_set    = u32(0x00020000)
	dependent_slice_segment_flag_set             = u32(0x00040000)
	slice_qp_delta                               = u32(0x00080000)
	different_slice_qp_delta                     = u32(0x00100000)
	max_enum_khr                                 = max_int
}
pub type VideoEncodeH265StdFlagsKHR = u32

pub enum VideoEncodeH265CtbSizeFlagBitsKHR as u32 {
	_16          = u32(0x00000001)
	_32          = u32(0x00000002)
	_64          = u32(0x00000004)
	max_enum_khr = max_int
}
pub type VideoEncodeH265CtbSizeFlagsKHR = u32

pub enum VideoEncodeH265TransformBlockSizeFlagBitsKHR as u32 {
	_4           = u32(0x00000001)
	_8           = u32(0x00000002)
	_16          = u32(0x00000004)
	_32          = u32(0x00000008)
	max_enum_khr = max_int
}
pub type VideoEncodeH265TransformBlockSizeFlagsKHR = u32

pub enum VideoEncodeH265RateControlFlagBitsKHR as u32 {
	attempt_hrd_compliance            = u32(0x00000001)
	regular_gop                       = u32(0x00000002)
	reference_pattern_flat            = u32(0x00000004)
	reference_pattern_dyadic          = u32(0x00000008)
	temporal_sub_layer_pattern_dyadic = u32(0x00000010)
	max_enum_khr                      = max_int
}
pub type VideoEncodeH265RateControlFlagsKHR = u32

// VideoEncodeH265CapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoEncodeH265CapabilitiesKHR = C.VkVideoEncodeH265CapabilitiesKHR

@[typedef]
pub struct C.VkVideoEncodeH265CapabilitiesKHR {
pub mut:
	sType                               StructureType = StructureType.video_encode_h265_capabilities_khr
	pNext                               voidptr       = unsafe { nil }
	flags                               VideoEncodeH265CapabilityFlagsKHR
	maxLevelIdc                         StdVideoH265LevelIdc
	maxSliceSegmentCount                u32
	maxTiles                            Extent2D
	ctbSizes                            VideoEncodeH265CtbSizeFlagsKHR
	transformBlockSizes                 VideoEncodeH265TransformBlockSizeFlagsKHR
	maxPPictureL0ReferenceCount         u32
	maxBPictureL0ReferenceCount         u32
	maxL1ReferenceCount                 u32
	maxSubLayerCount                    u32
	expectDyadicTemporalSubLayerPattern Bool32
	minQp                               i32
	maxQp                               i32
	prefersGopRemainingFrames           Bool32
	requiresGopRemainingFrames          Bool32
	stdSyntaxFlags                      VideoEncodeH265StdFlagsKHR
}

// VideoEncodeH265SessionCreateInfoKHR extends VkVideoSessionCreateInfoKHR
pub type VideoEncodeH265SessionCreateInfoKHR = C.VkVideoEncodeH265SessionCreateInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265SessionCreateInfoKHR {
pub mut:
	sType          StructureType = StructureType.video_encode_h265_session_create_info_khr
	pNext          voidptr       = unsafe { nil }
	useMaxLevelIdc Bool32
	maxLevelIdc    StdVideoH265LevelIdc
}

pub type VideoEncodeH265QpKHR = C.VkVideoEncodeH265QpKHR

@[typedef]
pub struct C.VkVideoEncodeH265QpKHR {
pub mut:
	qpI i32
	qpP i32
	qpB i32
}

// VideoEncodeH265QualityLevelPropertiesKHR extends VkVideoEncodeQualityLevelPropertiesKHR
pub type VideoEncodeH265QualityLevelPropertiesKHR = C.VkVideoEncodeH265QualityLevelPropertiesKHR

@[typedef]
pub struct C.VkVideoEncodeH265QualityLevelPropertiesKHR {
pub mut:
	sType                           StructureType = StructureType.video_encode_h265_quality_level_properties_khr
	pNext                           voidptr       = unsafe { nil }
	preferredRateControlFlags       VideoEncodeH265RateControlFlagsKHR
	preferredGopFrameCount          u32
	preferredIdrPeriod              u32
	preferredConsecutiveBFrameCount u32
	preferredSubLayerCount          u32
	preferredConstantQp             VideoEncodeH265QpKHR
	preferredMaxL0ReferenceCount    u32
	preferredMaxL1ReferenceCount    u32
}

// VideoEncodeH265SessionParametersAddInfoKHR extends VkVideoSessionParametersUpdateInfoKHR
pub type VideoEncodeH265SessionParametersAddInfoKHR = C.VkVideoEncodeH265SessionParametersAddInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265SessionParametersAddInfoKHR {
pub mut:
	sType       StructureType = StructureType.video_encode_h265_session_parameters_add_info_khr
	pNext       voidptr       = unsafe { nil }
	stdVPSCount u32
	pStdVPSs    &StdVideoH265VideoParameterSet
	stdSPSCount u32
	pStdSPSs    &StdVideoH265SequenceParameterSet
	stdPPSCount u32
	pStdPPSs    &StdVideoH265PictureParameterSet
}

// VideoEncodeH265SessionParametersCreateInfoKHR extends VkVideoSessionParametersCreateInfoKHR
pub type VideoEncodeH265SessionParametersCreateInfoKHR = C.VkVideoEncodeH265SessionParametersCreateInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265SessionParametersCreateInfoKHR {
pub mut:
	sType              StructureType = StructureType.video_encode_h265_session_parameters_create_info_khr
	pNext              voidptr       = unsafe { nil }
	maxStdVPSCount     u32
	maxStdSPSCount     u32
	maxStdPPSCount     u32
	pParametersAddInfo &VideoEncodeH265SessionParametersAddInfoKHR
}

// VideoEncodeH265SessionParametersGetInfoKHR extends VkVideoEncodeSessionParametersGetInfoKHR
pub type VideoEncodeH265SessionParametersGetInfoKHR = C.VkVideoEncodeH265SessionParametersGetInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265SessionParametersGetInfoKHR {
pub mut:
	sType       StructureType = StructureType.video_encode_h265_session_parameters_get_info_khr
	pNext       voidptr       = unsafe { nil }
	writeStdVPS Bool32
	writeStdSPS Bool32
	writeStdPPS Bool32
	stdVPSId    u32
	stdSPSId    u32
	stdPPSId    u32
}

// VideoEncodeH265SessionParametersFeedbackInfoKHR extends VkVideoEncodeSessionParametersFeedbackInfoKHR
pub type VideoEncodeH265SessionParametersFeedbackInfoKHR = C.VkVideoEncodeH265SessionParametersFeedbackInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265SessionParametersFeedbackInfoKHR {
pub mut:
	sType              StructureType = StructureType.video_encode_h265_session_parameters_feedback_info_khr
	pNext              voidptr       = unsafe { nil }
	hasStdVPSOverrides Bool32
	hasStdSPSOverrides Bool32
	hasStdPPSOverrides Bool32
}

pub type VideoEncodeH265NaluSliceSegmentInfoKHR = C.VkVideoEncodeH265NaluSliceSegmentInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265NaluSliceSegmentInfoKHR {
pub mut:
	sType                  StructureType = StructureType.video_encode_h265_nalu_slice_segment_info_khr
	pNext                  voidptr       = unsafe { nil }
	constantQp             i32
	pStdSliceSegmentHeader &StdVideoEncodeH265SliceSegmentHeader
}

// VideoEncodeH265PictureInfoKHR extends VkVideoEncodeInfoKHR
pub type VideoEncodeH265PictureInfoKHR = C.VkVideoEncodeH265PictureInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265PictureInfoKHR {
pub mut:
	sType                      StructureType = StructureType.video_encode_h265_picture_info_khr
	pNext                      voidptr       = unsafe { nil }
	naluSliceSegmentEntryCount u32
	pNaluSliceSegmentEntries   &VideoEncodeH265NaluSliceSegmentInfoKHR
	pStdPictureInfo            &StdVideoEncodeH265PictureInfo
}

// VideoEncodeH265DpbSlotInfoKHR extends VkVideoReferenceSlotInfoKHR
pub type VideoEncodeH265DpbSlotInfoKHR = C.VkVideoEncodeH265DpbSlotInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265DpbSlotInfoKHR {
pub mut:
	sType             StructureType = StructureType.video_encode_h265_dpb_slot_info_khr
	pNext             voidptr       = unsafe { nil }
	pStdReferenceInfo &StdVideoEncodeH265ReferenceInfo
}

// VideoEncodeH265ProfileInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub type VideoEncodeH265ProfileInfoKHR = C.VkVideoEncodeH265ProfileInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265ProfileInfoKHR {
pub mut:
	sType         StructureType = StructureType.video_encode_h265_profile_info_khr
	pNext         voidptr       = unsafe { nil }
	stdProfileIdc StdVideoH265ProfileIdc
}

// VideoEncodeH265RateControlInfoKHR extends VkVideoCodingControlInfoKHR,VkVideoBeginCodingInfoKHR
pub type VideoEncodeH265RateControlInfoKHR = C.VkVideoEncodeH265RateControlInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265RateControlInfoKHR {
pub mut:
	sType                  StructureType = StructureType.video_encode_h265_rate_control_info_khr
	pNext                  voidptr       = unsafe { nil }
	flags                  VideoEncodeH265RateControlFlagsKHR
	gopFrameCount          u32
	idrPeriod              u32
	consecutiveBFrameCount u32
	subLayerCount          u32
}

pub type VideoEncodeH265FrameSizeKHR = C.VkVideoEncodeH265FrameSizeKHR

@[typedef]
pub struct C.VkVideoEncodeH265FrameSizeKHR {
pub mut:
	frameISize u32
	framePSize u32
	frameBSize u32
}

// VideoEncodeH265RateControlLayerInfoKHR extends VkVideoEncodeRateControlLayerInfoKHR
pub type VideoEncodeH265RateControlLayerInfoKHR = C.VkVideoEncodeH265RateControlLayerInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265RateControlLayerInfoKHR {
pub mut:
	sType           StructureType = StructureType.video_encode_h265_rate_control_layer_info_khr
	pNext           voidptr       = unsafe { nil }
	useMinQp        Bool32
	minQp           VideoEncodeH265QpKHR
	useMaxQp        Bool32
	maxQp           VideoEncodeH265QpKHR
	useMaxFrameSize Bool32
	maxFrameSize    VideoEncodeH265FrameSizeKHR
}

// VideoEncodeH265GopRemainingFrameInfoKHR extends VkVideoBeginCodingInfoKHR
pub type VideoEncodeH265GopRemainingFrameInfoKHR = C.VkVideoEncodeH265GopRemainingFrameInfoKHR

@[typedef]
pub struct C.VkVideoEncodeH265GopRemainingFrameInfoKHR {
pub mut:
	sType                 StructureType = StructureType.video_encode_h265_gop_remaining_frame_info_khr
	pNext                 voidptr       = unsafe { nil }
	useGopRemainingFrames Bool32
	gopRemainingI         u32
	gopRemainingP         u32
	gopRemainingB         u32
}

pub const khr_video_decode_h264_spec_version = 9
pub const khr_video_decode_h264_extension_name = c'VK_KHR_video_decode_h264'

pub enum VideoDecodeH264PictureLayoutFlagBitsKHR as u32 {
	progressive                  = 0
	interlaced_interleaved_lines = u32(0x00000001)
	interlaced_separate_planes   = u32(0x00000002)
	max_enum_khr                 = max_int
}
pub type VideoDecodeH264PictureLayoutFlagsKHR = u32

// VideoDecodeH264ProfileInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub type VideoDecodeH264ProfileInfoKHR = C.VkVideoDecodeH264ProfileInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH264ProfileInfoKHR {
pub mut:
	sType         StructureType = StructureType.video_decode_h264_profile_info_khr
	pNext         voidptr       = unsafe { nil }
	stdProfileIdc StdVideoH264ProfileIdc
	pictureLayout VideoDecodeH264PictureLayoutFlagBitsKHR
}

// VideoDecodeH264CapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoDecodeH264CapabilitiesKHR = C.VkVideoDecodeH264CapabilitiesKHR

@[typedef]
pub struct C.VkVideoDecodeH264CapabilitiesKHR {
pub mut:
	sType                  StructureType = StructureType.video_decode_h264_capabilities_khr
	pNext                  voidptr       = unsafe { nil }
	maxLevelIdc            StdVideoH264LevelIdc
	fieldOffsetGranularity Offset2D
}

// VideoDecodeH264SessionParametersAddInfoKHR extends VkVideoSessionParametersUpdateInfoKHR
pub type VideoDecodeH264SessionParametersAddInfoKHR = C.VkVideoDecodeH264SessionParametersAddInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH264SessionParametersAddInfoKHR {
pub mut:
	sType       StructureType = StructureType.video_decode_h264_session_parameters_add_info_khr
	pNext       voidptr       = unsafe { nil }
	stdSPSCount u32
	pStdSPSs    &StdVideoH264SequenceParameterSet
	stdPPSCount u32
	pStdPPSs    &StdVideoH264PictureParameterSet
}

// VideoDecodeH264SessionParametersCreateInfoKHR extends VkVideoSessionParametersCreateInfoKHR
pub type VideoDecodeH264SessionParametersCreateInfoKHR = C.VkVideoDecodeH264SessionParametersCreateInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH264SessionParametersCreateInfoKHR {
pub mut:
	sType              StructureType = StructureType.video_decode_h264_session_parameters_create_info_khr
	pNext              voidptr       = unsafe { nil }
	maxStdSPSCount     u32
	maxStdPPSCount     u32
	pParametersAddInfo &VideoDecodeH264SessionParametersAddInfoKHR
}

// VideoDecodeH264PictureInfoKHR extends VkVideoDecodeInfoKHR
pub type VideoDecodeH264PictureInfoKHR = C.VkVideoDecodeH264PictureInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH264PictureInfoKHR {
pub mut:
	sType           StructureType = StructureType.video_decode_h264_picture_info_khr
	pNext           voidptr       = unsafe { nil }
	pStdPictureInfo &StdVideoDecodeH264PictureInfo
	sliceCount      u32
	pSliceOffsets   &u32
}

// VideoDecodeH264DpbSlotInfoKHR extends VkVideoReferenceSlotInfoKHR
pub type VideoDecodeH264DpbSlotInfoKHR = C.VkVideoDecodeH264DpbSlotInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH264DpbSlotInfoKHR {
pub mut:
	sType             StructureType = StructureType.video_decode_h264_dpb_slot_info_khr
	pNext             voidptr       = unsafe { nil }
	pStdReferenceInfo &StdVideoDecodeH264ReferenceInfo
}

pub const khr_dynamic_rendering_spec_version = 1
pub const khr_dynamic_rendering_extension_name = c'VK_KHR_dynamic_rendering'

pub type RenderingFlagsKHR = u32
pub type RenderingFlagBitsKHR = RenderingFlagBits

pub type RenderingInfoKHR = C.VkRenderingInfo

pub type RenderingAttachmentInfoKHR = C.VkRenderingAttachmentInfo

pub type PipelineRenderingCreateInfoKHR = C.VkPipelineRenderingCreateInfo

pub type PhysicalDeviceDynamicRenderingFeaturesKHR = C.VkPhysicalDeviceDynamicRenderingFeatures

pub type CommandBufferInheritanceRenderingInfoKHR = C.VkCommandBufferInheritanceRenderingInfo

@[keep_args_alive]
fn C.vkCmdBeginRenderingKHR(command_buffer CommandBuffer, p_rendering_info &RenderingInfo)

pub type PFN_vkCmdBeginRenderingKHR = fn (command_buffer CommandBuffer, p_rendering_info &RenderingInfo)

@[inline]
pub fn cmd_begin_rendering_khr(command_buffer CommandBuffer,
	p_rendering_info &RenderingInfo) {
	C.vkCmdBeginRenderingKHR(command_buffer, p_rendering_info)
}

@[keep_args_alive]
fn C.vkCmdEndRenderingKHR(command_buffer CommandBuffer)

pub type PFN_vkCmdEndRenderingKHR = fn (command_buffer CommandBuffer)

@[inline]
pub fn cmd_end_rendering_khr(command_buffer CommandBuffer) {
	C.vkCmdEndRenderingKHR(command_buffer)
}

pub const khr_multiview_spec_version = 1
pub const khr_multiview_extension_name = c'VK_KHR_multiview'

pub type RenderPassMultiviewCreateInfoKHR = C.VkRenderPassMultiviewCreateInfo

pub type PhysicalDeviceMultiviewFeaturesKHR = C.VkPhysicalDeviceMultiviewFeatures

pub type PhysicalDeviceMultiviewPropertiesKHR = C.VkPhysicalDeviceMultiviewProperties

pub const khr_get_physical_device_properties_2_spec_version = 2
pub const khr_get_physical_device_properties_2_extension_name = c'VK_KHR_get_physical_device_properties2'

pub type PhysicalDeviceFeatures2KHR = C.VkPhysicalDeviceFeatures2

pub type PhysicalDeviceProperties2KHR = C.VkPhysicalDeviceProperties2

pub type FormatProperties2KHR = C.VkFormatProperties2

pub type ImageFormatProperties2KHR = C.VkImageFormatProperties2

pub type PhysicalDeviceImageFormatInfo2KHR = C.VkPhysicalDeviceImageFormatInfo2

pub type QueueFamilyProperties2KHR = C.VkQueueFamilyProperties2

pub type PhysicalDeviceMemoryProperties2KHR = C.VkPhysicalDeviceMemoryProperties2

pub type SparseImageFormatProperties2KHR = C.VkSparseImageFormatProperties2

pub type PhysicalDeviceSparseImageFormatInfo2KHR = C.VkPhysicalDeviceSparseImageFormatInfo2

@[keep_args_alive]
fn C.vkGetPhysicalDeviceFeatures2KHR(physical_device PhysicalDevice, mut p_features PhysicalDeviceFeatures2)

pub type PFN_vkGetPhysicalDeviceFeatures2KHR = fn (physical_device PhysicalDevice, mut p_features PhysicalDeviceFeatures2)

@[inline]
pub fn get_physical_device_features2_khr(physical_device PhysicalDevice,
	mut p_features PhysicalDeviceFeatures2) {
	C.vkGetPhysicalDeviceFeatures2KHR(physical_device, mut p_features)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceProperties2KHR(physical_device PhysicalDevice, mut p_properties PhysicalDeviceProperties2)

pub type PFN_vkGetPhysicalDeviceProperties2KHR = fn (physical_device PhysicalDevice, mut p_properties PhysicalDeviceProperties2)

@[inline]
pub fn get_physical_device_properties2_khr(physical_device PhysicalDevice,
	mut p_properties PhysicalDeviceProperties2) {
	C.vkGetPhysicalDeviceProperties2KHR(physical_device, mut p_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceFormatProperties2KHR(physical_device PhysicalDevice, format Format, mut p_format_properties FormatProperties2)

pub type PFN_vkGetPhysicalDeviceFormatProperties2KHR = fn (physical_device PhysicalDevice, format Format, mut p_format_properties FormatProperties2)

@[inline]
pub fn get_physical_device_format_properties2_khr(physical_device PhysicalDevice,
	format Format,
	mut p_format_properties FormatProperties2) {
	C.vkGetPhysicalDeviceFormatProperties2KHR(physical_device, format, mut p_format_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceImageFormatProperties2KHR(physical_device PhysicalDevice, p_image_format_info &PhysicalDeviceImageFormatInfo2, mut p_image_format_properties ImageFormatProperties2) Result

pub type PFN_vkGetPhysicalDeviceImageFormatProperties2KHR = fn (physical_device PhysicalDevice, p_image_format_info &PhysicalDeviceImageFormatInfo2, mut p_image_format_properties ImageFormatProperties2) Result

@[inline]
pub fn get_physical_device_image_format_properties2_khr(physical_device PhysicalDevice,
	p_image_format_info &PhysicalDeviceImageFormatInfo2,
	mut p_image_format_properties ImageFormatProperties2) Result {
	return C.vkGetPhysicalDeviceImageFormatProperties2KHR(physical_device, p_image_format_info, mut
		p_image_format_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceQueueFamilyProperties2KHR(physical_device PhysicalDevice, p_queue_family_property_count &u32, mut p_queue_family_properties QueueFamilyProperties2)

pub type PFN_vkGetPhysicalDeviceQueueFamilyProperties2KHR = fn (physical_device PhysicalDevice, p_queue_family_property_count &u32, mut p_queue_family_properties QueueFamilyProperties2)

@[inline]
pub fn get_physical_device_queue_family_properties2_khr(physical_device PhysicalDevice,
	p_queue_family_property_count &u32,
	mut p_queue_family_properties QueueFamilyProperties2) {
	C.vkGetPhysicalDeviceQueueFamilyProperties2KHR(physical_device, p_queue_family_property_count, mut
		p_queue_family_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceMemoryProperties2KHR(physical_device PhysicalDevice, mut p_memory_properties PhysicalDeviceMemoryProperties2)

pub type PFN_vkGetPhysicalDeviceMemoryProperties2KHR = fn (physical_device PhysicalDevice, mut p_memory_properties PhysicalDeviceMemoryProperties2)

@[inline]
pub fn get_physical_device_memory_properties2_khr(physical_device PhysicalDevice,
	mut p_memory_properties PhysicalDeviceMemoryProperties2) {
	C.vkGetPhysicalDeviceMemoryProperties2KHR(physical_device, mut p_memory_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceSparseImageFormatProperties2KHR(physical_device PhysicalDevice, p_format_info &PhysicalDeviceSparseImageFormatInfo2, p_property_count &u32, mut p_properties SparseImageFormatProperties2)

pub type PFN_vkGetPhysicalDeviceSparseImageFormatProperties2KHR = fn (physical_device PhysicalDevice, p_format_info &PhysicalDeviceSparseImageFormatInfo2, p_property_count &u32, mut p_properties SparseImageFormatProperties2)

@[inline]
pub fn get_physical_device_sparse_image_format_properties2_khr(physical_device PhysicalDevice,
	p_format_info &PhysicalDeviceSparseImageFormatInfo2,
	p_property_count &u32,
	mut p_properties SparseImageFormatProperties2) {
	C.vkGetPhysicalDeviceSparseImageFormatProperties2KHR(physical_device, p_format_info,
		p_property_count, mut p_properties)
}

pub const khr_device_group_spec_version = 4
pub const khr_device_group_extension_name = c'VK_KHR_device_group'

pub type PeerMemoryFeatureFlagsKHR = u32
pub type PeerMemoryFeatureFlagBitsKHR = PeerMemoryFeatureFlagBits

pub type MemoryAllocateFlagsKHR = u32
pub type MemoryAllocateFlagBitsKHR = MemoryAllocateFlagBits

pub type MemoryAllocateFlagsInfoKHR = C.VkMemoryAllocateFlagsInfo

pub type DeviceGroupRenderPassBeginInfoKHR = C.VkDeviceGroupRenderPassBeginInfo

pub type DeviceGroupCommandBufferBeginInfoKHR = C.VkDeviceGroupCommandBufferBeginInfo

pub type DeviceGroupSubmitInfoKHR = C.VkDeviceGroupSubmitInfo

pub type DeviceGroupBindSparseInfoKHR = C.VkDeviceGroupBindSparseInfo

pub type BindBufferMemoryDeviceGroupInfoKHR = C.VkBindBufferMemoryDeviceGroupInfo

pub type BindImageMemoryDeviceGroupInfoKHR = C.VkBindImageMemoryDeviceGroupInfo

@[keep_args_alive]
fn C.vkGetDeviceGroupPeerMemoryFeaturesKHR(device Device, heap_index u32, local_device_index u32, remote_device_index u32, p_peer_memory_features &PeerMemoryFeatureFlags)

pub type PFN_vkGetDeviceGroupPeerMemoryFeaturesKHR = fn (device Device, heap_index u32, local_device_index u32, remote_device_index u32, p_peer_memory_features &PeerMemoryFeatureFlags)

@[inline]
pub fn get_device_group_peer_memory_features_khr(device Device,
	heap_index u32,
	local_device_index u32,
	remote_device_index u32,
	p_peer_memory_features &PeerMemoryFeatureFlags) {
	C.vkGetDeviceGroupPeerMemoryFeaturesKHR(device, heap_index, local_device_index, remote_device_index,
		p_peer_memory_features)
}

@[keep_args_alive]
fn C.vkCmdSetDeviceMaskKHR(command_buffer CommandBuffer, device_mask u32)

pub type PFN_vkCmdSetDeviceMaskKHR = fn (command_buffer CommandBuffer, device_mask u32)

@[inline]
pub fn cmd_set_device_mask_khr(command_buffer CommandBuffer,
	device_mask u32) {
	C.vkCmdSetDeviceMaskKHR(command_buffer, device_mask)
}

@[keep_args_alive]
fn C.vkCmdDispatchBaseKHR(command_buffer CommandBuffer, base_group_x u32, base_group_y u32, base_group_z u32, group_count_x u32, group_count_y u32, group_count_z u32)

pub type PFN_vkCmdDispatchBaseKHR = fn (command_buffer CommandBuffer, base_group_x u32, base_group_y u32, base_group_z u32, group_count_x u32, group_count_y u32, group_count_z u32)

@[inline]
pub fn cmd_dispatch_base_khr(command_buffer CommandBuffer,
	base_group_x u32,
	base_group_y u32,
	base_group_z u32,
	group_count_x u32,
	group_count_y u32,
	group_count_z u32) {
	C.vkCmdDispatchBaseKHR(command_buffer, base_group_x, base_group_y, base_group_z, group_count_x,
		group_count_y, group_count_z)
}

pub const khr_shader_draw_parameters_spec_version = 1
pub const khr_shader_draw_parameters_extension_name = c'VK_KHR_shader_draw_parameters'

pub const khr_maintenance_1_spec_version = 2
pub const khr_maintenance_1_extension_name = c'VK_KHR_maintenance1'
// VK_KHR_MAINTENANCE1_SPEC_VERSION is a deprecated alias
pub const khr_maintenance1_spec_version = khr_maintenance_1_spec_version
// VK_KHR_MAINTENANCE1_EXTENSION_NAME is a deprecated alias
pub const khr_maintenance1_extension_name = khr_maintenance_1_extension_name

pub type CommandPoolTrimFlagsKHR = u32

@[keep_args_alive]
fn C.vkTrimCommandPoolKHR(device Device, command_pool CommandPool, flags CommandPoolTrimFlags)

pub type PFN_vkTrimCommandPoolKHR = fn (device Device, command_pool CommandPool, flags CommandPoolTrimFlags)

@[inline]
pub fn trim_command_pool_khr(device Device,
	command_pool CommandPool,
	flags CommandPoolTrimFlags) {
	C.vkTrimCommandPoolKHR(device, command_pool, flags)
}

pub const khr_device_group_creation_spec_version = 1
pub const khr_device_group_creation_extension_name = c'VK_KHR_device_group_creation'
pub const max_device_group_size_khr = max_device_group_size

pub type PhysicalDeviceGroupPropertiesKHR = C.VkPhysicalDeviceGroupProperties

pub type DeviceGroupDeviceCreateInfoKHR = C.VkDeviceGroupDeviceCreateInfo

@[keep_args_alive]
fn C.vkEnumeratePhysicalDeviceGroupsKHR(instance Instance, p_physical_device_group_count &u32, mut p_physical_device_group_properties PhysicalDeviceGroupProperties) Result

pub type PFN_vkEnumeratePhysicalDeviceGroupsKHR = fn (instance Instance, p_physical_device_group_count &u32, mut p_physical_device_group_properties PhysicalDeviceGroupProperties) Result

@[inline]
pub fn enumerate_physical_device_groups_khr(instance Instance,
	p_physical_device_group_count &u32,
	mut p_physical_device_group_properties PhysicalDeviceGroupProperties) Result {
	return C.vkEnumeratePhysicalDeviceGroupsKHR(instance, p_physical_device_group_count, mut
		p_physical_device_group_properties)
}

pub const khr_external_memory_capabilities_spec_version = 1
pub const khr_external_memory_capabilities_extension_name = c'VK_KHR_external_memory_capabilities'
pub const luid_size_khr = luid_size

pub type ExternalMemoryHandleTypeFlagsKHR = u32
pub type ExternalMemoryHandleTypeFlagBitsKHR = ExternalMemoryHandleTypeFlagBits

pub type ExternalMemoryFeatureFlagsKHR = u32
pub type ExternalMemoryFeatureFlagBitsKHR = ExternalMemoryFeatureFlagBits

pub type ExternalMemoryPropertiesKHR = C.VkExternalMemoryProperties

pub type PhysicalDeviceExternalImageFormatInfoKHR = C.VkPhysicalDeviceExternalImageFormatInfo

pub type ExternalImageFormatPropertiesKHR = C.VkExternalImageFormatProperties

pub type PhysicalDeviceExternalBufferInfoKHR = C.VkPhysicalDeviceExternalBufferInfo

pub type ExternalBufferPropertiesKHR = C.VkExternalBufferProperties

pub type PhysicalDeviceIDPropertiesKHR = C.VkPhysicalDeviceIDProperties

@[keep_args_alive]
fn C.vkGetPhysicalDeviceExternalBufferPropertiesKHR(physical_device PhysicalDevice, p_external_buffer_info &PhysicalDeviceExternalBufferInfo, mut p_external_buffer_properties ExternalBufferProperties)

pub type PFN_vkGetPhysicalDeviceExternalBufferPropertiesKHR = fn (physical_device PhysicalDevice, p_external_buffer_info &PhysicalDeviceExternalBufferInfo, mut p_external_buffer_properties ExternalBufferProperties)

@[inline]
pub fn get_physical_device_external_buffer_properties_khr(physical_device PhysicalDevice,
	p_external_buffer_info &PhysicalDeviceExternalBufferInfo,
	mut p_external_buffer_properties ExternalBufferProperties) {
	C.vkGetPhysicalDeviceExternalBufferPropertiesKHR(physical_device, p_external_buffer_info, mut
		p_external_buffer_properties)
}

pub const khr_external_memory_spec_version = 1
pub const khr_external_memory_extension_name = c'VK_KHR_external_memory'
pub const queue_family_external_khr = queue_family_external

pub type ExternalMemoryImageCreateInfoKHR = C.VkExternalMemoryImageCreateInfo

pub type ExternalMemoryBufferCreateInfoKHR = C.VkExternalMemoryBufferCreateInfo

pub type ExportMemoryAllocateInfoKHR = C.VkExportMemoryAllocateInfo

pub const khr_external_memory_fd_spec_version = 1
pub const khr_external_memory_fd_extension_name = c'VK_KHR_external_memory_fd'
// ImportMemoryFdInfoKHR extends VkMemoryAllocateInfo
pub type ImportMemoryFdInfoKHR = C.VkImportMemoryFdInfoKHR

@[typedef]
pub struct C.VkImportMemoryFdInfoKHR {
pub mut:
	sType      StructureType = StructureType.import_memory_fd_info_khr
	pNext      voidptr       = unsafe { nil }
	handleType ExternalMemoryHandleTypeFlagBits
	fd         int
}

pub type MemoryFdPropertiesKHR = C.VkMemoryFdPropertiesKHR

@[typedef]
pub struct C.VkMemoryFdPropertiesKHR {
pub mut:
	sType          StructureType = StructureType.memory_fd_properties_khr
	pNext          voidptr       = unsafe { nil }
	memoryTypeBits u32
}

pub type MemoryGetFdInfoKHR = C.VkMemoryGetFdInfoKHR

@[typedef]
pub struct C.VkMemoryGetFdInfoKHR {
pub mut:
	sType      StructureType = StructureType.memory_get_fd_info_khr
	pNext      voidptr       = unsafe { nil }
	memory     DeviceMemory
	handleType ExternalMemoryHandleTypeFlagBits
}

@[keep_args_alive]
fn C.vkGetMemoryFdKHR(device Device, p_get_fd_info &MemoryGetFdInfoKHR, p_fd &int) Result

pub type PFN_vkGetMemoryFdKHR = fn (device Device, p_get_fd_info &MemoryGetFdInfoKHR, p_fd &int) Result

@[inline]
pub fn get_memory_fd_khr(device Device,
	p_get_fd_info &MemoryGetFdInfoKHR,
	p_fd &int) Result {
	return C.vkGetMemoryFdKHR(device, p_get_fd_info, p_fd)
}

@[keep_args_alive]
fn C.vkGetMemoryFdPropertiesKHR(device Device, handle_type ExternalMemoryHandleTypeFlagBits, fd int, mut p_memory_fd_properties MemoryFdPropertiesKHR) Result

pub type PFN_vkGetMemoryFdPropertiesKHR = fn (device Device, handle_type ExternalMemoryHandleTypeFlagBits, fd int, mut p_memory_fd_properties MemoryFdPropertiesKHR) Result

@[inline]
pub fn get_memory_fd_properties_khr(device Device,
	handle_type ExternalMemoryHandleTypeFlagBits,
	fd int,
	mut p_memory_fd_properties MemoryFdPropertiesKHR) Result {
	return C.vkGetMemoryFdPropertiesKHR(device, handle_type, fd, mut p_memory_fd_properties)
}

pub const khr_external_semaphore_capabilities_spec_version = 1
pub const khr_external_semaphore_capabilities_extension_name = c'VK_KHR_external_semaphore_capabilities'

pub type ExternalSemaphoreHandleTypeFlagsKHR = u32
pub type ExternalSemaphoreHandleTypeFlagBitsKHR = ExternalSemaphoreHandleTypeFlagBits

pub type ExternalSemaphoreFeatureFlagsKHR = u32
pub type ExternalSemaphoreFeatureFlagBitsKHR = ExternalSemaphoreFeatureFlagBits

pub type PhysicalDeviceExternalSemaphoreInfoKHR = C.VkPhysicalDeviceExternalSemaphoreInfo

pub type ExternalSemaphorePropertiesKHR = C.VkExternalSemaphoreProperties

@[keep_args_alive]
fn C.vkGetPhysicalDeviceExternalSemaphorePropertiesKHR(physical_device PhysicalDevice, p_external_semaphore_info &PhysicalDeviceExternalSemaphoreInfo, mut p_external_semaphore_properties ExternalSemaphoreProperties)

pub type PFN_vkGetPhysicalDeviceExternalSemaphorePropertiesKHR = fn (physical_device PhysicalDevice, p_external_semaphore_info &PhysicalDeviceExternalSemaphoreInfo, mut p_external_semaphore_properties ExternalSemaphoreProperties)

@[inline]
pub fn get_physical_device_external_semaphore_properties_khr(physical_device PhysicalDevice,
	p_external_semaphore_info &PhysicalDeviceExternalSemaphoreInfo,
	mut p_external_semaphore_properties ExternalSemaphoreProperties) {
	C.vkGetPhysicalDeviceExternalSemaphorePropertiesKHR(physical_device, p_external_semaphore_info, mut
		p_external_semaphore_properties)
}

pub const khr_external_semaphore_spec_version = 1
pub const khr_external_semaphore_extension_name = c'VK_KHR_external_semaphore'

pub type SemaphoreImportFlagsKHR = u32
pub type SemaphoreImportFlagBitsKHR = SemaphoreImportFlagBits

pub type ExportSemaphoreCreateInfoKHR = C.VkExportSemaphoreCreateInfo

pub const khr_external_semaphore_fd_spec_version = 1
pub const khr_external_semaphore_fd_extension_name = c'VK_KHR_external_semaphore_fd'

pub type ImportSemaphoreFdInfoKHR = C.VkImportSemaphoreFdInfoKHR

@[typedef]
pub struct C.VkImportSemaphoreFdInfoKHR {
pub mut:
	sType      StructureType = StructureType.import_semaphore_fd_info_khr
	pNext      voidptr       = unsafe { nil }
	semaphore  Semaphore
	flags      SemaphoreImportFlags
	handleType ExternalSemaphoreHandleTypeFlagBits
	fd         int
}

pub type SemaphoreGetFdInfoKHR = C.VkSemaphoreGetFdInfoKHR

@[typedef]
pub struct C.VkSemaphoreGetFdInfoKHR {
pub mut:
	sType      StructureType = StructureType.semaphore_get_fd_info_khr
	pNext      voidptr       = unsafe { nil }
	semaphore  Semaphore
	handleType ExternalSemaphoreHandleTypeFlagBits
}

@[keep_args_alive]
fn C.vkImportSemaphoreFdKHR(device Device, p_import_semaphore_fd_info &ImportSemaphoreFdInfoKHR) Result

pub type PFN_vkImportSemaphoreFdKHR = fn (device Device, p_import_semaphore_fd_info &ImportSemaphoreFdInfoKHR) Result

@[inline]
pub fn import_semaphore_fd_khr(device Device,
	p_import_semaphore_fd_info &ImportSemaphoreFdInfoKHR) Result {
	return C.vkImportSemaphoreFdKHR(device, p_import_semaphore_fd_info)
}

@[keep_args_alive]
fn C.vkGetSemaphoreFdKHR(device Device, p_get_fd_info &SemaphoreGetFdInfoKHR, p_fd &int) Result

pub type PFN_vkGetSemaphoreFdKHR = fn (device Device, p_get_fd_info &SemaphoreGetFdInfoKHR, p_fd &int) Result

@[inline]
pub fn get_semaphore_fd_khr(device Device,
	p_get_fd_info &SemaphoreGetFdInfoKHR,
	p_fd &int) Result {
	return C.vkGetSemaphoreFdKHR(device, p_get_fd_info, p_fd)
}

pub const khr_push_descriptor_spec_version = 2
pub const khr_push_descriptor_extension_name = c'VK_KHR_push_descriptor'

pub type PhysicalDevicePushDescriptorPropertiesKHR = C.VkPhysicalDevicePushDescriptorProperties

@[keep_args_alive]
fn C.vkCmdPushDescriptorSetKHR(command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, layout PipelineLayout, set u32, descriptor_write_count u32, p_descriptor_writes &WriteDescriptorSet)

pub type PFN_vkCmdPushDescriptorSetKHR = fn (command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, layout PipelineLayout, set u32, descriptor_write_count u32, p_descriptor_writes &WriteDescriptorSet)

@[inline]
pub fn cmd_push_descriptor_set_khr(command_buffer CommandBuffer,
	pipeline_bind_point PipelineBindPoint,
	layout PipelineLayout,
	set u32,
	descriptor_write_count u32,
	p_descriptor_writes &WriteDescriptorSet) {
	C.vkCmdPushDescriptorSetKHR(command_buffer, pipeline_bind_point, layout, set, descriptor_write_count,
		p_descriptor_writes)
}

@[keep_args_alive]
fn C.vkCmdPushDescriptorSetWithTemplateKHR(command_buffer CommandBuffer, descriptor_update_template DescriptorUpdateTemplate, layout PipelineLayout, set u32, p_data voidptr)

pub type PFN_vkCmdPushDescriptorSetWithTemplateKHR = fn (command_buffer CommandBuffer, descriptor_update_template DescriptorUpdateTemplate, layout PipelineLayout, set u32, p_data voidptr)

@[inline]
pub fn cmd_push_descriptor_set_with_template_khr(command_buffer CommandBuffer,
	descriptor_update_template DescriptorUpdateTemplate,
	layout PipelineLayout,
	set u32,
	p_data voidptr) {
	C.vkCmdPushDescriptorSetWithTemplateKHR(command_buffer, descriptor_update_template,
		layout, set, p_data)
}

pub const khr_shader_float16_int8_spec_version = 1
pub const khr_shader_float16_int8_extension_name = c'VK_KHR_shader_float16_int8'

pub type PhysicalDeviceShaderFloat16Int8FeaturesKHR = C.VkPhysicalDeviceShaderFloat16Int8Features

pub type PhysicalDeviceFloat16Int8FeaturesKHR = C.VkPhysicalDeviceShaderFloat16Int8Features

pub const khr_16bit_storage_spec_version = 1
pub const khr_16bit_storage_extension_name = c'VK_KHR_16bit_storage'

pub type PhysicalDevice16BitStorageFeaturesKHR = C.VkPhysicalDevice16BitStorageFeatures

pub const khr_incremental_present_spec_version = 2
pub const khr_incremental_present_extension_name = c'VK_KHR_incremental_present'

pub type RectLayerKHR = C.VkRectLayerKHR

@[typedef]
pub struct C.VkRectLayerKHR {
pub mut:
	offset Offset2D
	extent Extent2D
	layer  u32
}

pub type PresentRegionKHR = C.VkPresentRegionKHR

@[typedef]
pub struct C.VkPresentRegionKHR {
pub mut:
	rectangleCount u32
	pRectangles    &RectLayerKHR
}

// PresentRegionsKHR extends VkPresentInfoKHR
pub type PresentRegionsKHR = C.VkPresentRegionsKHR

@[typedef]
pub struct C.VkPresentRegionsKHR {
pub mut:
	sType          StructureType = StructureType.present_regions_khr
	pNext          voidptr       = unsafe { nil }
	swapchainCount u32
	pRegions       &PresentRegionKHR
}

pub type DescriptorUpdateTemplateKHR = voidptr

pub const khr_descriptor_update_template_spec_version = 1
pub const khr_descriptor_update_template_extension_name = c'VK_KHR_descriptor_update_template'

pub type DescriptorUpdateTemplateTypeKHR = DescriptorUpdateTemplateType

pub type DescriptorUpdateTemplateCreateFlagsKHR = u32
pub type DescriptorUpdateTemplateEntryKHR = C.VkDescriptorUpdateTemplateEntry

pub type DescriptorUpdateTemplateCreateInfoKHR = C.VkDescriptorUpdateTemplateCreateInfo

@[keep_args_alive]
fn C.vkCreateDescriptorUpdateTemplateKHR(device Device, p_create_info &DescriptorUpdateTemplateCreateInfo, p_allocator &AllocationCallbacks, p_descriptor_update_template &DescriptorUpdateTemplate) Result

pub type PFN_vkCreateDescriptorUpdateTemplateKHR = fn (device Device, p_create_info &DescriptorUpdateTemplateCreateInfo, p_allocator &AllocationCallbacks, p_descriptor_update_template &DescriptorUpdateTemplate) Result

@[inline]
pub fn create_descriptor_update_template_khr(device Device,
	p_create_info &DescriptorUpdateTemplateCreateInfo,
	p_allocator &AllocationCallbacks,
	p_descriptor_update_template &DescriptorUpdateTemplate) Result {
	return C.vkCreateDescriptorUpdateTemplateKHR(device, p_create_info, p_allocator, p_descriptor_update_template)
}

@[keep_args_alive]
fn C.vkDestroyDescriptorUpdateTemplateKHR(device Device, descriptor_update_template DescriptorUpdateTemplate, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyDescriptorUpdateTemplateKHR = fn (device Device, descriptor_update_template DescriptorUpdateTemplate, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_descriptor_update_template_khr(device Device,
	descriptor_update_template DescriptorUpdateTemplate,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyDescriptorUpdateTemplateKHR(device, descriptor_update_template, p_allocator)
}

@[keep_args_alive]
fn C.vkUpdateDescriptorSetWithTemplateKHR(device Device, descriptor_set DescriptorSet, descriptor_update_template DescriptorUpdateTemplate, p_data voidptr)

pub type PFN_vkUpdateDescriptorSetWithTemplateKHR = fn (device Device, descriptor_set DescriptorSet, descriptor_update_template DescriptorUpdateTemplate, p_data voidptr)

@[inline]
pub fn update_descriptor_set_with_template_khr(device Device,
	descriptor_set DescriptorSet,
	descriptor_update_template DescriptorUpdateTemplate,
	p_data voidptr) {
	C.vkUpdateDescriptorSetWithTemplateKHR(device, descriptor_set, descriptor_update_template,
		p_data)
}

pub const khr_imageless_framebuffer_spec_version = 1
pub const khr_imageless_framebuffer_extension_name = c'VK_KHR_imageless_framebuffer'

pub type PhysicalDeviceImagelessFramebufferFeaturesKHR = C.VkPhysicalDeviceImagelessFramebufferFeatures

pub type FramebufferAttachmentsCreateInfoKHR = C.VkFramebufferAttachmentsCreateInfo

pub type FramebufferAttachmentImageInfoKHR = C.VkFramebufferAttachmentImageInfo

pub type RenderPassAttachmentBeginInfoKHR = C.VkRenderPassAttachmentBeginInfo

pub const khr_create_renderpass_2_spec_version = 1
pub const khr_create_renderpass_2_extension_name = c'VK_KHR_create_renderpass2'

pub type RenderPassCreateInfo2KHR = C.VkRenderPassCreateInfo2

pub type AttachmentDescription2KHR = C.VkAttachmentDescription2

pub type AttachmentReference2KHR = C.VkAttachmentReference2

pub type SubpassDescription2KHR = C.VkSubpassDescription2

pub type SubpassDependency2KHR = C.VkSubpassDependency2

pub type SubpassBeginInfoKHR = C.VkSubpassBeginInfo

pub type SubpassEndInfoKHR = C.VkSubpassEndInfo

@[keep_args_alive]
fn C.vkCreateRenderPass2KHR(device Device, p_create_info &RenderPassCreateInfo2, p_allocator &AllocationCallbacks, p_render_pass &RenderPass) Result

pub type PFN_vkCreateRenderPass2KHR = fn (device Device, p_create_info &RenderPassCreateInfo2, p_allocator &AllocationCallbacks, p_render_pass &RenderPass) Result

@[inline]
pub fn create_render_pass2_khr(device Device,
	p_create_info &RenderPassCreateInfo2,
	p_allocator &AllocationCallbacks,
	p_render_pass &RenderPass) Result {
	return C.vkCreateRenderPass2KHR(device, p_create_info, p_allocator, p_render_pass)
}

@[keep_args_alive]
fn C.vkCmdBeginRenderPass2KHR(command_buffer CommandBuffer, p_render_pass_begin &RenderPassBeginInfo, p_subpass_begin_info &SubpassBeginInfo)

pub type PFN_vkCmdBeginRenderPass2KHR = fn (command_buffer CommandBuffer, p_render_pass_begin &RenderPassBeginInfo, p_subpass_begin_info &SubpassBeginInfo)

@[inline]
pub fn cmd_begin_render_pass2_khr(command_buffer CommandBuffer,
	p_render_pass_begin &RenderPassBeginInfo,
	p_subpass_begin_info &SubpassBeginInfo) {
	C.vkCmdBeginRenderPass2KHR(command_buffer, p_render_pass_begin, p_subpass_begin_info)
}

@[keep_args_alive]
fn C.vkCmdNextSubpass2KHR(command_buffer CommandBuffer, p_subpass_begin_info &SubpassBeginInfo, p_subpass_end_info &SubpassEndInfo)

pub type PFN_vkCmdNextSubpass2KHR = fn (command_buffer CommandBuffer, p_subpass_begin_info &SubpassBeginInfo, p_subpass_end_info &SubpassEndInfo)

@[inline]
pub fn cmd_next_subpass2_khr(command_buffer CommandBuffer,
	p_subpass_begin_info &SubpassBeginInfo,
	p_subpass_end_info &SubpassEndInfo) {
	C.vkCmdNextSubpass2KHR(command_buffer, p_subpass_begin_info, p_subpass_end_info)
}

@[keep_args_alive]
fn C.vkCmdEndRenderPass2KHR(command_buffer CommandBuffer, p_subpass_end_info &SubpassEndInfo)

pub type PFN_vkCmdEndRenderPass2KHR = fn (command_buffer CommandBuffer, p_subpass_end_info &SubpassEndInfo)

@[inline]
pub fn cmd_end_render_pass2_khr(command_buffer CommandBuffer,
	p_subpass_end_info &SubpassEndInfo) {
	C.vkCmdEndRenderPass2KHR(command_buffer, p_subpass_end_info)
}

pub const khr_shared_presentable_image_spec_version = 1
pub const khr_shared_presentable_image_extension_name = c'VK_KHR_shared_presentable_image'
// SharedPresentSurfaceCapabilitiesKHR extends VkSurfaceCapabilities2KHR
pub type SharedPresentSurfaceCapabilitiesKHR = C.VkSharedPresentSurfaceCapabilitiesKHR

@[typedef]
pub struct C.VkSharedPresentSurfaceCapabilitiesKHR {
pub mut:
	sType                            StructureType = StructureType.shared_present_surface_capabilities_khr
	pNext                            voidptr       = unsafe { nil }
	sharedPresentSupportedUsageFlags ImageUsageFlags
}

@[keep_args_alive]
fn C.vkGetSwapchainStatusKHR(device Device, swapchain SwapchainKHR) Result

pub type PFN_vkGetSwapchainStatusKHR = fn (device Device, swapchain SwapchainKHR) Result

@[inline]
pub fn get_swapchain_status_khr(device Device,
	swapchain SwapchainKHR) Result {
	return C.vkGetSwapchainStatusKHR(device, swapchain)
}

pub const khr_external_fence_capabilities_spec_version = 1
pub const khr_external_fence_capabilities_extension_name = c'VK_KHR_external_fence_capabilities'

pub type ExternalFenceHandleTypeFlagsKHR = u32
pub type ExternalFenceHandleTypeFlagBitsKHR = ExternalFenceHandleTypeFlagBits

pub type ExternalFenceFeatureFlagsKHR = u32
pub type ExternalFenceFeatureFlagBitsKHR = ExternalFenceFeatureFlagBits

pub type PhysicalDeviceExternalFenceInfoKHR = C.VkPhysicalDeviceExternalFenceInfo

pub type ExternalFencePropertiesKHR = C.VkExternalFenceProperties

@[keep_args_alive]
fn C.vkGetPhysicalDeviceExternalFencePropertiesKHR(physical_device PhysicalDevice, p_external_fence_info &PhysicalDeviceExternalFenceInfo, mut p_external_fence_properties ExternalFenceProperties)

pub type PFN_vkGetPhysicalDeviceExternalFencePropertiesKHR = fn (physical_device PhysicalDevice, p_external_fence_info &PhysicalDeviceExternalFenceInfo, mut p_external_fence_properties ExternalFenceProperties)

@[inline]
pub fn get_physical_device_external_fence_properties_khr(physical_device PhysicalDevice,
	p_external_fence_info &PhysicalDeviceExternalFenceInfo,
	mut p_external_fence_properties ExternalFenceProperties) {
	C.vkGetPhysicalDeviceExternalFencePropertiesKHR(physical_device, p_external_fence_info, mut
		p_external_fence_properties)
}

pub const khr_external_fence_spec_version = 1
pub const khr_external_fence_extension_name = c'VK_KHR_external_fence'

pub type FenceImportFlagsKHR = u32
pub type FenceImportFlagBitsKHR = FenceImportFlagBits

pub type ExportFenceCreateInfoKHR = C.VkExportFenceCreateInfo

pub const khr_external_fence_fd_spec_version = 1
pub const khr_external_fence_fd_extension_name = c'VK_KHR_external_fence_fd'

pub type ImportFenceFdInfoKHR = C.VkImportFenceFdInfoKHR

@[typedef]
pub struct C.VkImportFenceFdInfoKHR {
pub mut:
	sType      StructureType = StructureType.import_fence_fd_info_khr
	pNext      voidptr       = unsafe { nil }
	fence      Fence
	flags      FenceImportFlags
	handleType ExternalFenceHandleTypeFlagBits
	fd         int
}

pub type FenceGetFdInfoKHR = C.VkFenceGetFdInfoKHR

@[typedef]
pub struct C.VkFenceGetFdInfoKHR {
pub mut:
	sType      StructureType = StructureType.fence_get_fd_info_khr
	pNext      voidptr       = unsafe { nil }
	fence      Fence
	handleType ExternalFenceHandleTypeFlagBits
}

@[keep_args_alive]
fn C.vkImportFenceFdKHR(device Device, p_import_fence_fd_info &ImportFenceFdInfoKHR) Result

pub type PFN_vkImportFenceFdKHR = fn (device Device, p_import_fence_fd_info &ImportFenceFdInfoKHR) Result

@[inline]
pub fn import_fence_fd_khr(device Device,
	p_import_fence_fd_info &ImportFenceFdInfoKHR) Result {
	return C.vkImportFenceFdKHR(device, p_import_fence_fd_info)
}

@[keep_args_alive]
fn C.vkGetFenceFdKHR(device Device, p_get_fd_info &FenceGetFdInfoKHR, p_fd &int) Result

pub type PFN_vkGetFenceFdKHR = fn (device Device, p_get_fd_info &FenceGetFdInfoKHR, p_fd &int) Result

@[inline]
pub fn get_fence_fd_khr(device Device,
	p_get_fd_info &FenceGetFdInfoKHR,
	p_fd &int) Result {
	return C.vkGetFenceFdKHR(device, p_get_fd_info, p_fd)
}

pub const khr_performance_query_spec_version = 1
pub const khr_performance_query_extension_name = c'VK_KHR_performance_query'

pub enum PerformanceCounterUnitKHR as u32 {
	generic          = 0
	percentage       = 1
	nanoseconds      = 2
	bytes            = 3
	bytes_per_second = 4
	kelvin           = 5
	watts            = 6
	volts            = 7
	amps             = 8
	hertz            = 9
	cycles           = 10
	max_enum_khr     = max_int
}

pub enum PerformanceCounterScopeKHR as u32 {
	command_buffer = 0
	render_pass    = 1
	command        = 2
	max_enum_khr   = max_int
}

pub enum PerformanceCounterStorageKHR as u32 {
	int32        = 0
	int64        = 1
	uint32       = 2
	uint64       = 3
	float32      = 4
	float64      = 5
	max_enum_khr = max_int
}

pub enum PerformanceCounterDescriptionFlagBitsKHR as u32 {
	performance_impacting = u32(0x00000001)
	concurrently_impacted = u32(0x00000002)
	max_enum_khr          = max_int
}
pub type PerformanceCounterDescriptionFlagsKHR = u32

pub enum AcquireProfilingLockFlagBitsKHR as u32 {
	max_enum_khr = max_int
}
pub type AcquireProfilingLockFlagsKHR = u32

// PhysicalDevicePerformanceQueryFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePerformanceQueryFeaturesKHR = C.VkPhysicalDevicePerformanceQueryFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDevicePerformanceQueryFeaturesKHR {
pub mut:
	sType                                StructureType = StructureType.physical_device_performance_query_features_khr
	pNext                                voidptr       = unsafe { nil }
	performanceCounterQueryPools         Bool32
	performanceCounterMultipleQueryPools Bool32
}

// PhysicalDevicePerformanceQueryPropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDevicePerformanceQueryPropertiesKHR = C.VkPhysicalDevicePerformanceQueryPropertiesKHR

@[typedef]
pub struct C.VkPhysicalDevicePerformanceQueryPropertiesKHR {
pub mut:
	sType                         StructureType = StructureType.physical_device_performance_query_properties_khr
	pNext                         voidptr       = unsafe { nil }
	allowCommandBufferQueryCopies Bool32
}

pub type PerformanceCounterKHR = C.VkPerformanceCounterKHR

@[typedef]
pub struct C.VkPerformanceCounterKHR {
pub mut:
	sType   StructureType = StructureType.performance_counter_khr
	pNext   voidptr       = unsafe { nil }
	unit    PerformanceCounterUnitKHR
	scope   PerformanceCounterScopeKHR
	storage PerformanceCounterStorageKHR
	uuid    [uuid_size]u8
}

pub type PerformanceCounterDescriptionKHR = C.VkPerformanceCounterDescriptionKHR

@[typedef]
pub struct C.VkPerformanceCounterDescriptionKHR {
pub mut:
	sType       StructureType = StructureType.performance_counter_description_khr
	pNext       voidptr       = unsafe { nil }
	flags       PerformanceCounterDescriptionFlagsKHR
	name        [max_description_size]char
	category    [max_description_size]char
	description [max_description_size]char
}

// QueryPoolPerformanceCreateInfoKHR extends VkQueryPoolCreateInfo
pub type QueryPoolPerformanceCreateInfoKHR = C.VkQueryPoolPerformanceCreateInfoKHR

@[typedef]
pub struct C.VkQueryPoolPerformanceCreateInfoKHR {
pub mut:
	sType             StructureType = StructureType.query_pool_performance_create_info_khr
	pNext             voidptr       = unsafe { nil }
	queueFamilyIndex  u32
	counterIndexCount u32
	pCounterIndices   &u32
}

pub type PerformanceCounterResultKHR = C.VkPerformanceCounterResultKHR

@[typedef]
pub union C.VkPerformanceCounterResultKHR {
pub mut:
	int32   i32
	int64   i64
	uint32  u32
	uint64  u64
	float32 f32
	float64 f64
}

pub type AcquireProfilingLockInfoKHR = C.VkAcquireProfilingLockInfoKHR

@[typedef]
pub struct C.VkAcquireProfilingLockInfoKHR {
pub mut:
	sType   StructureType = StructureType.acquire_profiling_lock_info_khr
	pNext   voidptr       = unsafe { nil }
	flags   AcquireProfilingLockFlagsKHR
	timeout u64
}

// PerformanceQuerySubmitInfoKHR extends VkSubmitInfo,VkSubmitInfo2
pub type PerformanceQuerySubmitInfoKHR = C.VkPerformanceQuerySubmitInfoKHR

@[typedef]
pub struct C.VkPerformanceQuerySubmitInfoKHR {
pub mut:
	sType            StructureType = StructureType.performance_query_submit_info_khr
	pNext            voidptr       = unsafe { nil }
	counterPassIndex u32
}

@[keep_args_alive]
fn C.vkEnumeratePhysicalDeviceQueueFamilyPerformanceQueryCountersKHR(physical_device PhysicalDevice, queue_family_index u32, p_counter_count &u32, mut p_counters PerformanceCounterKHR, mut p_counter_descriptions PerformanceCounterDescriptionKHR) Result

pub type PFN_vkEnumeratePhysicalDeviceQueueFamilyPerformanceQueryCountersKHR = fn (physical_device PhysicalDevice, queue_family_index u32, p_counter_count &u32, mut p_counters PerformanceCounterKHR, mut p_counter_descriptions PerformanceCounterDescriptionKHR) Result

@[inline]
pub fn enumerate_physical_device_queue_family_performance_query_counters_khr(physical_device PhysicalDevice,
	queue_family_index u32,
	p_counter_count &u32,
	mut p_counters PerformanceCounterKHR,
	mut p_counter_descriptions PerformanceCounterDescriptionKHR) Result {
	return C.vkEnumeratePhysicalDeviceQueueFamilyPerformanceQueryCountersKHR(physical_device,
		queue_family_index, p_counter_count, mut p_counters, mut p_counter_descriptions)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceQueueFamilyPerformanceQueryPassesKHR(physical_device PhysicalDevice, p_performance_query_create_info &QueryPoolPerformanceCreateInfoKHR, p_num_passes &u32)

pub type PFN_vkGetPhysicalDeviceQueueFamilyPerformanceQueryPassesKHR = fn (physical_device PhysicalDevice, p_performance_query_create_info &QueryPoolPerformanceCreateInfoKHR, p_num_passes &u32)

@[inline]
pub fn get_physical_device_queue_family_performance_query_passes_khr(physical_device PhysicalDevice,
	p_performance_query_create_info &QueryPoolPerformanceCreateInfoKHR,
	p_num_passes &u32) {
	C.vkGetPhysicalDeviceQueueFamilyPerformanceQueryPassesKHR(physical_device, p_performance_query_create_info,
		p_num_passes)
}

@[keep_args_alive]
fn C.vkAcquireProfilingLockKHR(device Device, p_info &AcquireProfilingLockInfoKHR) Result

pub type PFN_vkAcquireProfilingLockKHR = fn (device Device, p_info &AcquireProfilingLockInfoKHR) Result

@[inline]
pub fn acquire_profiling_lock_khr(device Device,
	p_info &AcquireProfilingLockInfoKHR) Result {
	return C.vkAcquireProfilingLockKHR(device, p_info)
}

@[keep_args_alive]
fn C.vkReleaseProfilingLockKHR(device Device)

pub type PFN_vkReleaseProfilingLockKHR = fn (device Device)

@[inline]
pub fn release_profiling_lock_khr(device Device) {
	C.vkReleaseProfilingLockKHR(device)
}

pub const khr_maintenance_2_spec_version = 1
pub const khr_maintenance_2_extension_name = c'VK_KHR_maintenance2'
// VK_KHR_MAINTENANCE2_SPEC_VERSION is a deprecated alias
pub const khr_maintenance2_spec_version = khr_maintenance_2_spec_version
// VK_KHR_MAINTENANCE2_EXTENSION_NAME is a deprecated alias
pub const khr_maintenance2_extension_name = khr_maintenance_2_extension_name

pub type PointClippingBehaviorKHR = PointClippingBehavior

pub type TessellationDomainOriginKHR = TessellationDomainOrigin

pub type PhysicalDevicePointClippingPropertiesKHR = C.VkPhysicalDevicePointClippingProperties

pub type RenderPassInputAttachmentAspectCreateInfoKHR = C.VkRenderPassInputAttachmentAspectCreateInfo

pub type InputAttachmentAspectReferenceKHR = C.VkInputAttachmentAspectReference

pub type ImageViewUsageCreateInfoKHR = C.VkImageViewUsageCreateInfo

pub type PipelineTessellationDomainOriginStateCreateInfoKHR = C.VkPipelineTessellationDomainOriginStateCreateInfo

pub const khr_get_surface_capabilities_2_spec_version = 1
pub const khr_get_surface_capabilities_2_extension_name = c'VK_KHR_get_surface_capabilities2'

pub type PhysicalDeviceSurfaceInfo2KHR = C.VkPhysicalDeviceSurfaceInfo2KHR

@[typedef]
pub struct C.VkPhysicalDeviceSurfaceInfo2KHR {
pub mut:
	sType   StructureType = StructureType.physical_device_surface_info2_khr
	pNext   voidptr       = unsafe { nil }
	surface SurfaceKHR
}

pub type SurfaceCapabilities2KHR = C.VkSurfaceCapabilities2KHR

@[typedef]
pub struct C.VkSurfaceCapabilities2KHR {
pub mut:
	sType               StructureType = StructureType.surface_capabilities2_khr
	pNext               voidptr       = unsafe { nil }
	surfaceCapabilities SurfaceCapabilitiesKHR
}

pub type SurfaceFormat2KHR = C.VkSurfaceFormat2KHR

@[typedef]
pub struct C.VkSurfaceFormat2KHR {
pub mut:
	sType         StructureType = StructureType.surface_format2_khr
	pNext         voidptr       = unsafe { nil }
	surfaceFormat SurfaceFormatKHR
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceSurfaceCapabilities2KHR(physical_device PhysicalDevice, p_surface_info &PhysicalDeviceSurfaceInfo2KHR, mut p_surface_capabilities SurfaceCapabilities2KHR) Result

pub type PFN_vkGetPhysicalDeviceSurfaceCapabilities2KHR = fn (physical_device PhysicalDevice, p_surface_info &PhysicalDeviceSurfaceInfo2KHR, mut p_surface_capabilities SurfaceCapabilities2KHR) Result

@[inline]
pub fn get_physical_device_surface_capabilities2_khr(physical_device PhysicalDevice,
	p_surface_info &PhysicalDeviceSurfaceInfo2KHR,
	mut p_surface_capabilities SurfaceCapabilities2KHR) Result {
	return C.vkGetPhysicalDeviceSurfaceCapabilities2KHR(physical_device, p_surface_info, mut
		p_surface_capabilities)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceSurfaceFormats2KHR(physical_device PhysicalDevice, p_surface_info &PhysicalDeviceSurfaceInfo2KHR, p_surface_format_count &u32, mut p_surface_formats SurfaceFormat2KHR) Result

pub type PFN_vkGetPhysicalDeviceSurfaceFormats2KHR = fn (physical_device PhysicalDevice, p_surface_info &PhysicalDeviceSurfaceInfo2KHR, p_surface_format_count &u32, mut p_surface_formats SurfaceFormat2KHR) Result

@[inline]
pub fn get_physical_device_surface_formats2_khr(physical_device PhysicalDevice,
	p_surface_info &PhysicalDeviceSurfaceInfo2KHR,
	p_surface_format_count &u32,
	mut p_surface_formats SurfaceFormat2KHR) Result {
	return C.vkGetPhysicalDeviceSurfaceFormats2KHR(physical_device, p_surface_info, p_surface_format_count, mut
		p_surface_formats)
}

pub const khr_variable_pointers_spec_version = 1
pub const khr_variable_pointers_extension_name = c'VK_KHR_variable_pointers'

pub type PhysicalDeviceVariablePointerFeaturesKHR = C.VkPhysicalDeviceVariablePointersFeatures

pub type PhysicalDeviceVariablePointersFeaturesKHR = C.VkPhysicalDeviceVariablePointersFeatures

pub const khr_get_display_properties_2_spec_version = 1
pub const khr_get_display_properties_2_extension_name = c'VK_KHR_get_display_properties2'

pub type DisplayProperties2KHR = C.VkDisplayProperties2KHR

@[typedef]
pub struct C.VkDisplayProperties2KHR {
pub mut:
	sType             StructureType = StructureType.display_properties2_khr
	pNext             voidptr       = unsafe { nil }
	displayProperties DisplayPropertiesKHR
}

pub type DisplayPlaneProperties2KHR = C.VkDisplayPlaneProperties2KHR

@[typedef]
pub struct C.VkDisplayPlaneProperties2KHR {
pub mut:
	sType                  StructureType = StructureType.display_plane_properties2_khr
	pNext                  voidptr       = unsafe { nil }
	displayPlaneProperties DisplayPlanePropertiesKHR
}

pub type DisplayModeProperties2KHR = C.VkDisplayModeProperties2KHR

@[typedef]
pub struct C.VkDisplayModeProperties2KHR {
pub mut:
	sType                 StructureType = StructureType.display_mode_properties2_khr
	pNext                 voidptr       = unsafe { nil }
	displayModeProperties DisplayModePropertiesKHR
}

pub type DisplayPlaneInfo2KHR = C.VkDisplayPlaneInfo2KHR

@[typedef]
pub struct C.VkDisplayPlaneInfo2KHR {
pub mut:
	sType      StructureType = StructureType.display_plane_info2_khr
	pNext      voidptr       = unsafe { nil }
	mode       DisplayModeKHR
	planeIndex u32
}

pub type DisplayPlaneCapabilities2KHR = C.VkDisplayPlaneCapabilities2KHR

@[typedef]
pub struct C.VkDisplayPlaneCapabilities2KHR {
pub mut:
	sType        StructureType = StructureType.display_plane_capabilities2_khr
	pNext        voidptr       = unsafe { nil }
	capabilities DisplayPlaneCapabilitiesKHR
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceDisplayProperties2KHR(physical_device PhysicalDevice, p_property_count &u32, mut p_properties DisplayProperties2KHR) Result

pub type PFN_vkGetPhysicalDeviceDisplayProperties2KHR = fn (physical_device PhysicalDevice, p_property_count &u32, mut p_properties DisplayProperties2KHR) Result

@[inline]
pub fn get_physical_device_display_properties2_khr(physical_device PhysicalDevice,
	p_property_count &u32,
	mut p_properties DisplayProperties2KHR) Result {
	return C.vkGetPhysicalDeviceDisplayProperties2KHR(physical_device, p_property_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceDisplayPlaneProperties2KHR(physical_device PhysicalDevice, p_property_count &u32, mut p_properties DisplayPlaneProperties2KHR) Result

pub type PFN_vkGetPhysicalDeviceDisplayPlaneProperties2KHR = fn (physical_device PhysicalDevice, p_property_count &u32, mut p_properties DisplayPlaneProperties2KHR) Result

@[inline]
pub fn get_physical_device_display_plane_properties2_khr(physical_device PhysicalDevice,
	p_property_count &u32,
	mut p_properties DisplayPlaneProperties2KHR) Result {
	return C.vkGetPhysicalDeviceDisplayPlaneProperties2KHR(physical_device, p_property_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkGetDisplayModeProperties2KHR(physical_device PhysicalDevice, display DisplayKHR, p_property_count &u32, mut p_properties DisplayModeProperties2KHR) Result

pub type PFN_vkGetDisplayModeProperties2KHR = fn (physical_device PhysicalDevice, display DisplayKHR, p_property_count &u32, mut p_properties DisplayModeProperties2KHR) Result

@[inline]
pub fn get_display_mode_properties2_khr(physical_device PhysicalDevice,
	display DisplayKHR,
	p_property_count &u32,
	mut p_properties DisplayModeProperties2KHR) Result {
	return C.vkGetDisplayModeProperties2KHR(physical_device, display, p_property_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkGetDisplayPlaneCapabilities2KHR(physical_device PhysicalDevice, p_display_plane_info &DisplayPlaneInfo2KHR, mut p_capabilities DisplayPlaneCapabilities2KHR) Result

pub type PFN_vkGetDisplayPlaneCapabilities2KHR = fn (physical_device PhysicalDevice, p_display_plane_info &DisplayPlaneInfo2KHR, mut p_capabilities DisplayPlaneCapabilities2KHR) Result

@[inline]
pub fn get_display_plane_capabilities2_khr(physical_device PhysicalDevice,
	p_display_plane_info &DisplayPlaneInfo2KHR,
	mut p_capabilities DisplayPlaneCapabilities2KHR) Result {
	return C.vkGetDisplayPlaneCapabilities2KHR(physical_device, p_display_plane_info, mut
		p_capabilities)
}

pub const khr_dedicated_allocation_spec_version = 3
pub const khr_dedicated_allocation_extension_name = c'VK_KHR_dedicated_allocation'

pub type MemoryDedicatedRequirementsKHR = C.VkMemoryDedicatedRequirements

pub type MemoryDedicatedAllocateInfoKHR = C.VkMemoryDedicatedAllocateInfo

pub const khr_storage_buffer_storage_class_spec_version = 1
pub const khr_storage_buffer_storage_class_extension_name = c'VK_KHR_storage_buffer_storage_class'

pub const khr_shader_bfloat16_spec_version = 1
pub const khr_shader_bfloat16_extension_name = c'VK_KHR_shader_bfloat16'
// PhysicalDeviceShaderBfloat16FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderBfloat16FeaturesKHR = C.VkPhysicalDeviceShaderBfloat16FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceShaderBfloat16FeaturesKHR {
pub mut:
	sType                           StructureType = StructureType.physical_device_shader_bfloat16_features_khr
	pNext                           voidptr       = unsafe { nil }
	shaderBFloat16Type              Bool32
	shaderBFloat16DotProduct        Bool32
	shaderBFloat16CooperativeMatrix Bool32
}

pub const khr_relaxed_block_layout_spec_version = 1
pub const khr_relaxed_block_layout_extension_name = c'VK_KHR_relaxed_block_layout'

pub const khr_get_memory_requirements_2_spec_version = 1
pub const khr_get_memory_requirements_2_extension_name = c'VK_KHR_get_memory_requirements2'

pub type BufferMemoryRequirementsInfo2KHR = C.VkBufferMemoryRequirementsInfo2

pub type ImageMemoryRequirementsInfo2KHR = C.VkImageMemoryRequirementsInfo2

pub type ImageSparseMemoryRequirementsInfo2KHR = C.VkImageSparseMemoryRequirementsInfo2

pub type MemoryRequirements2KHR = C.VkMemoryRequirements2

pub type SparseImageMemoryRequirements2KHR = C.VkSparseImageMemoryRequirements2

@[keep_args_alive]
fn C.vkGetImageMemoryRequirements2KHR(device Device, p_info &ImageMemoryRequirementsInfo2, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetImageMemoryRequirements2KHR = fn (device Device, p_info &ImageMemoryRequirementsInfo2, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_image_memory_requirements2_khr(device Device,
	p_info &ImageMemoryRequirementsInfo2,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetImageMemoryRequirements2KHR(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetBufferMemoryRequirements2KHR(device Device, p_info &BufferMemoryRequirementsInfo2, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetBufferMemoryRequirements2KHR = fn (device Device, p_info &BufferMemoryRequirementsInfo2, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_buffer_memory_requirements2_khr(device Device,
	p_info &BufferMemoryRequirementsInfo2,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetBufferMemoryRequirements2KHR(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetImageSparseMemoryRequirements2KHR(device Device, p_info &ImageSparseMemoryRequirementsInfo2, p_sparse_memory_requirement_count &u32, mut p_sparse_memory_requirements SparseImageMemoryRequirements2)

pub type PFN_vkGetImageSparseMemoryRequirements2KHR = fn (device Device, p_info &ImageSparseMemoryRequirementsInfo2, p_sparse_memory_requirement_count &u32, mut p_sparse_memory_requirements SparseImageMemoryRequirements2)

@[inline]
pub fn get_image_sparse_memory_requirements2_khr(device Device,
	p_info &ImageSparseMemoryRequirementsInfo2,
	p_sparse_memory_requirement_count &u32,
	mut p_sparse_memory_requirements SparseImageMemoryRequirements2) {
	C.vkGetImageSparseMemoryRequirements2KHR(device, p_info, p_sparse_memory_requirement_count, mut
		p_sparse_memory_requirements)
}

pub const khr_image_format_list_spec_version = 1
pub const khr_image_format_list_extension_name = c'VK_KHR_image_format_list'

pub type ImageFormatListCreateInfoKHR = C.VkImageFormatListCreateInfo

pub type SamplerYcbcrConversionKHR = voidptr

pub const khr_sampler_ycbcr_conversion_spec_version = 14
pub const khr_sampler_ycbcr_conversion_extension_name = c'VK_KHR_sampler_ycbcr_conversion'

pub type SamplerYcbcrModelConversionKHR = SamplerYcbcrModelConversion

pub type SamplerYcbcrRangeKHR = SamplerYcbcrRange

pub type ChromaLocationKHR = ChromaLocation

pub type SamplerYcbcrConversionCreateInfoKHR = C.VkSamplerYcbcrConversionCreateInfo

pub type SamplerYcbcrConversionInfoKHR = C.VkSamplerYcbcrConversionInfo

pub type BindImagePlaneMemoryInfoKHR = C.VkBindImagePlaneMemoryInfo

pub type ImagePlaneMemoryRequirementsInfoKHR = C.VkImagePlaneMemoryRequirementsInfo

pub type PhysicalDeviceSamplerYcbcrConversionFeaturesKHR = C.VkPhysicalDeviceSamplerYcbcrConversionFeatures

pub type SamplerYcbcrConversionImageFormatPropertiesKHR = C.VkSamplerYcbcrConversionImageFormatProperties

@[keep_args_alive]
fn C.vkCreateSamplerYcbcrConversionKHR(device Device, p_create_info &SamplerYcbcrConversionCreateInfo, p_allocator &AllocationCallbacks, p_ycbcr_conversion &SamplerYcbcrConversion) Result

pub type PFN_vkCreateSamplerYcbcrConversionKHR = fn (device Device, p_create_info &SamplerYcbcrConversionCreateInfo, p_allocator &AllocationCallbacks, p_ycbcr_conversion &SamplerYcbcrConversion) Result

@[inline]
pub fn create_sampler_ycbcr_conversion_khr(device Device,
	p_create_info &SamplerYcbcrConversionCreateInfo,
	p_allocator &AllocationCallbacks,
	p_ycbcr_conversion &SamplerYcbcrConversion) Result {
	return C.vkCreateSamplerYcbcrConversionKHR(device, p_create_info, p_allocator, p_ycbcr_conversion)
}

@[keep_args_alive]
fn C.vkDestroySamplerYcbcrConversionKHR(device Device, ycbcr_conversion SamplerYcbcrConversion, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroySamplerYcbcrConversionKHR = fn (device Device, ycbcr_conversion SamplerYcbcrConversion, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_sampler_ycbcr_conversion_khr(device Device,
	ycbcr_conversion SamplerYcbcrConversion,
	p_allocator &AllocationCallbacks) {
	C.vkDestroySamplerYcbcrConversionKHR(device, ycbcr_conversion, p_allocator)
}

pub const khr_bind_memory_2_spec_version = 1
pub const khr_bind_memory_2_extension_name = c'VK_KHR_bind_memory2'

pub type BindBufferMemoryInfoKHR = C.VkBindBufferMemoryInfo

pub type BindImageMemoryInfoKHR = C.VkBindImageMemoryInfo

@[keep_args_alive]
fn C.vkBindBufferMemory2KHR(device Device, bind_info_count u32, p_bind_infos &BindBufferMemoryInfo) Result

pub type PFN_vkBindBufferMemory2KHR = fn (device Device, bind_info_count u32, p_bind_infos &BindBufferMemoryInfo) Result

@[inline]
pub fn bind_buffer_memory2_khr(device Device,
	bind_info_count u32,
	p_bind_infos &BindBufferMemoryInfo) Result {
	return C.vkBindBufferMemory2KHR(device, bind_info_count, p_bind_infos)
}

@[keep_args_alive]
fn C.vkBindImageMemory2KHR(device Device, bind_info_count u32, p_bind_infos &BindImageMemoryInfo) Result

pub type PFN_vkBindImageMemory2KHR = fn (device Device, bind_info_count u32, p_bind_infos &BindImageMemoryInfo) Result

@[inline]
pub fn bind_image_memory2_khr(device Device,
	bind_info_count u32,
	p_bind_infos &BindImageMemoryInfo) Result {
	return C.vkBindImageMemory2KHR(device, bind_info_count, p_bind_infos)
}

pub const khr_maintenance_3_spec_version = 1
pub const khr_maintenance_3_extension_name = c'VK_KHR_maintenance3'
// VK_KHR_MAINTENANCE3_SPEC_VERSION is a deprecated alias
pub const khr_maintenance3_spec_version = khr_maintenance_3_spec_version
// VK_KHR_MAINTENANCE3_EXTENSION_NAME is a deprecated alias
pub const khr_maintenance3_extension_name = khr_maintenance_3_extension_name

pub type PhysicalDeviceMaintenance3PropertiesKHR = C.VkPhysicalDeviceMaintenance3Properties

pub type DescriptorSetLayoutSupportKHR = C.VkDescriptorSetLayoutSupport

@[keep_args_alive]
fn C.vkGetDescriptorSetLayoutSupportKHR(device Device, p_create_info &DescriptorSetLayoutCreateInfo, mut p_support DescriptorSetLayoutSupport)

pub type PFN_vkGetDescriptorSetLayoutSupportKHR = fn (device Device, p_create_info &DescriptorSetLayoutCreateInfo, mut p_support DescriptorSetLayoutSupport)

@[inline]
pub fn get_descriptor_set_layout_support_khr(device Device,
	p_create_info &DescriptorSetLayoutCreateInfo,
	mut p_support DescriptorSetLayoutSupport) {
	C.vkGetDescriptorSetLayoutSupportKHR(device, p_create_info, mut p_support)
}

pub const khr_draw_indirect_count_spec_version = 1
pub const khr_draw_indirect_count_extension_name = c'VK_KHR_draw_indirect_count'

@[keep_args_alive]
fn C.vkCmdDrawIndirectCountKHR(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

pub type PFN_vkCmdDrawIndirectCountKHR = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_indirect_count_khr(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	count_buffer Buffer,
	count_buffer_offset DeviceSize,
	max_draw_count u32,
	stride u32) {
	C.vkCmdDrawIndirectCountKHR(command_buffer, buffer, offset, count_buffer, count_buffer_offset,
		max_draw_count, stride)
}

@[keep_args_alive]
fn C.vkCmdDrawIndexedIndirectCountKHR(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

pub type PFN_vkCmdDrawIndexedIndirectCountKHR = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_indexed_indirect_count_khr(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	count_buffer Buffer,
	count_buffer_offset DeviceSize,
	max_draw_count u32,
	stride u32) {
	C.vkCmdDrawIndexedIndirectCountKHR(command_buffer, buffer, offset, count_buffer, count_buffer_offset,
		max_draw_count, stride)
}

pub const khr_shader_subgroup_extended_types_spec_version = 1
pub const khr_shader_subgroup_extended_types_extension_name = c'VK_KHR_shader_subgroup_extended_types'

pub type PhysicalDeviceShaderSubgroupExtendedTypesFeaturesKHR = C.VkPhysicalDeviceShaderSubgroupExtendedTypesFeatures

pub const khr_8bit_storage_spec_version = 1
pub const khr_8bit_storage_extension_name = c'VK_KHR_8bit_storage'

pub type PhysicalDevice8BitStorageFeaturesKHR = C.VkPhysicalDevice8BitStorageFeatures

pub const khr_shader_atomic_int64_spec_version = 1
pub const khr_shader_atomic_int64_extension_name = c'VK_KHR_shader_atomic_int64'

pub type PhysicalDeviceShaderAtomicInt64FeaturesKHR = C.VkPhysicalDeviceShaderAtomicInt64Features

pub const khr_shader_clock_spec_version = 1
pub const khr_shader_clock_extension_name = c'VK_KHR_shader_clock'
// PhysicalDeviceShaderClockFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderClockFeaturesKHR = C.VkPhysicalDeviceShaderClockFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceShaderClockFeaturesKHR {
pub mut:
	sType               StructureType = StructureType.physical_device_shader_clock_features_khr
	pNext               voidptr       = unsafe { nil }
	shaderSubgroupClock Bool32
	shaderDeviceClock   Bool32
}

pub const khr_video_decode_h265_spec_version = 8
pub const khr_video_decode_h265_extension_name = c'VK_KHR_video_decode_h265'
// VideoDecodeH265ProfileInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub type VideoDecodeH265ProfileInfoKHR = C.VkVideoDecodeH265ProfileInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH265ProfileInfoKHR {
pub mut:
	sType         StructureType = StructureType.video_decode_h265_profile_info_khr
	pNext         voidptr       = unsafe { nil }
	stdProfileIdc StdVideoH265ProfileIdc
}

// VideoDecodeH265CapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoDecodeH265CapabilitiesKHR = C.VkVideoDecodeH265CapabilitiesKHR

@[typedef]
pub struct C.VkVideoDecodeH265CapabilitiesKHR {
pub mut:
	sType       StructureType = StructureType.video_decode_h265_capabilities_khr
	pNext       voidptr       = unsafe { nil }
	maxLevelIdc StdVideoH265LevelIdc
}

// VideoDecodeH265SessionParametersAddInfoKHR extends VkVideoSessionParametersUpdateInfoKHR
pub type VideoDecodeH265SessionParametersAddInfoKHR = C.VkVideoDecodeH265SessionParametersAddInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH265SessionParametersAddInfoKHR {
pub mut:
	sType       StructureType = StructureType.video_decode_h265_session_parameters_add_info_khr
	pNext       voidptr       = unsafe { nil }
	stdVPSCount u32
	pStdVPSs    &StdVideoH265VideoParameterSet
	stdSPSCount u32
	pStdSPSs    &StdVideoH265SequenceParameterSet
	stdPPSCount u32
	pStdPPSs    &StdVideoH265PictureParameterSet
}

// VideoDecodeH265SessionParametersCreateInfoKHR extends VkVideoSessionParametersCreateInfoKHR
pub type VideoDecodeH265SessionParametersCreateInfoKHR = C.VkVideoDecodeH265SessionParametersCreateInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH265SessionParametersCreateInfoKHR {
pub mut:
	sType              StructureType = StructureType.video_decode_h265_session_parameters_create_info_khr
	pNext              voidptr       = unsafe { nil }
	maxStdVPSCount     u32
	maxStdSPSCount     u32
	maxStdPPSCount     u32
	pParametersAddInfo &VideoDecodeH265SessionParametersAddInfoKHR
}

// VideoDecodeH265PictureInfoKHR extends VkVideoDecodeInfoKHR
pub type VideoDecodeH265PictureInfoKHR = C.VkVideoDecodeH265PictureInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH265PictureInfoKHR {
pub mut:
	sType                StructureType = StructureType.video_decode_h265_picture_info_khr
	pNext                voidptr       = unsafe { nil }
	pStdPictureInfo      &StdVideoDecodeH265PictureInfo
	sliceSegmentCount    u32
	pSliceSegmentOffsets &u32
}

// VideoDecodeH265DpbSlotInfoKHR extends VkVideoReferenceSlotInfoKHR
pub type VideoDecodeH265DpbSlotInfoKHR = C.VkVideoDecodeH265DpbSlotInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH265DpbSlotInfoKHR {
pub mut:
	sType             StructureType = StructureType.video_decode_h265_dpb_slot_info_khr
	pNext             voidptr       = unsafe { nil }
	pStdReferenceInfo &StdVideoDecodeH265ReferenceInfo
}

pub const khr_global_priority_spec_version = 1
pub const khr_global_priority_extension_name = c'VK_KHR_global_priority'
pub const max_global_priority_size_khr = max_global_priority_size

pub type QueueGlobalPriorityKHR = QueueGlobalPriority

pub type DeviceQueueGlobalPriorityCreateInfoKHR = C.VkDeviceQueueGlobalPriorityCreateInfo

pub type PhysicalDeviceGlobalPriorityQueryFeaturesKHR = C.VkPhysicalDeviceGlobalPriorityQueryFeatures

pub type QueueFamilyGlobalPriorityPropertiesKHR = C.VkQueueFamilyGlobalPriorityProperties

pub const khr_driver_properties_spec_version = 1
pub const khr_driver_properties_extension_name = c'VK_KHR_driver_properties'
pub const max_driver_name_size_khr = max_driver_name_size
pub const max_driver_info_size_khr = max_driver_info_size

pub type DriverIdKHR = DriverId

pub type ConformanceVersionKHR = C.VkConformanceVersion

pub type PhysicalDeviceDriverPropertiesKHR = C.VkPhysicalDeviceDriverProperties

pub const khr_shader_float_controls_spec_version = 4
pub const khr_shader_float_controls_extension_name = c'VK_KHR_shader_float_controls'

pub type ShaderFloatControlsIndependenceKHR = ShaderFloatControlsIndependence

pub type PhysicalDeviceFloatControlsPropertiesKHR = C.VkPhysicalDeviceFloatControlsProperties

pub const khr_depth_stencil_resolve_spec_version = 1
pub const khr_depth_stencil_resolve_extension_name = c'VK_KHR_depth_stencil_resolve'

pub type ResolveModeFlagBitsKHR = ResolveModeFlagBits

pub type ResolveModeFlagsKHR = u32
pub type SubpassDescriptionDepthStencilResolveKHR = C.VkSubpassDescriptionDepthStencilResolve

pub type PhysicalDeviceDepthStencilResolvePropertiesKHR = C.VkPhysicalDeviceDepthStencilResolveProperties

pub const khr_swapchain_mutable_format_spec_version = 1
pub const khr_swapchain_mutable_format_extension_name = c'VK_KHR_swapchain_mutable_format'

pub const khr_timeline_semaphore_spec_version = 2
pub const khr_timeline_semaphore_extension_name = c'VK_KHR_timeline_semaphore'

pub type SemaphoreTypeKHR = SemaphoreType

pub type SemaphoreWaitFlagBitsKHR = SemaphoreWaitFlagBits

pub type SemaphoreWaitFlagsKHR = u32
pub type PhysicalDeviceTimelineSemaphoreFeaturesKHR = C.VkPhysicalDeviceTimelineSemaphoreFeatures

pub type PhysicalDeviceTimelineSemaphorePropertiesKHR = C.VkPhysicalDeviceTimelineSemaphoreProperties

pub type SemaphoreTypeCreateInfoKHR = C.VkSemaphoreTypeCreateInfo

pub type TimelineSemaphoreSubmitInfoKHR = C.VkTimelineSemaphoreSubmitInfo

pub type SemaphoreWaitInfoKHR = C.VkSemaphoreWaitInfo

pub type SemaphoreSignalInfoKHR = C.VkSemaphoreSignalInfo

@[keep_args_alive]
fn C.vkGetSemaphoreCounterValueKHR(device Device, semaphore Semaphore, p_value &u64) Result

pub type PFN_vkGetSemaphoreCounterValueKHR = fn (device Device, semaphore Semaphore, p_value &u64) Result

@[inline]
pub fn get_semaphore_counter_value_khr(device Device,
	semaphore Semaphore,
	p_value &u64) Result {
	return C.vkGetSemaphoreCounterValueKHR(device, semaphore, p_value)
}

@[keep_args_alive]
fn C.vkWaitSemaphoresKHR(device Device, p_wait_info &SemaphoreWaitInfo, timeout u64) Result

pub type PFN_vkWaitSemaphoresKHR = fn (device Device, p_wait_info &SemaphoreWaitInfo, timeout u64) Result

@[inline]
pub fn wait_semaphores_khr(device Device,
	p_wait_info &SemaphoreWaitInfo,
	timeout u64) Result {
	return C.vkWaitSemaphoresKHR(device, p_wait_info, timeout)
}

@[keep_args_alive]
fn C.vkSignalSemaphoreKHR(device Device, p_signal_info &SemaphoreSignalInfo) Result

pub type PFN_vkSignalSemaphoreKHR = fn (device Device, p_signal_info &SemaphoreSignalInfo) Result

@[inline]
pub fn signal_semaphore_khr(device Device,
	p_signal_info &SemaphoreSignalInfo) Result {
	return C.vkSignalSemaphoreKHR(device, p_signal_info)
}

pub const khr_vulkan_memory_model_spec_version = 3
pub const khr_vulkan_memory_model_extension_name = c'VK_KHR_vulkan_memory_model'

pub type PhysicalDeviceVulkanMemoryModelFeaturesKHR = C.VkPhysicalDeviceVulkanMemoryModelFeatures

pub const khr_shader_terminate_invocation_spec_version = 1
pub const khr_shader_terminate_invocation_extension_name = c'VK_KHR_shader_terminate_invocation'

pub type PhysicalDeviceShaderTerminateInvocationFeaturesKHR = C.VkPhysicalDeviceShaderTerminateInvocationFeatures

pub const khr_fragment_shading_rate_spec_version = 2
pub const khr_fragment_shading_rate_extension_name = c'VK_KHR_fragment_shading_rate'

pub enum FragmentShadingRateCombinerOpKHR as u32 {
	keep         = 0
	replace      = 1
	min          = 2
	max          = 3
	mul          = 4
	max_enum_khr = max_int
}
// FragmentShadingRateAttachmentInfoKHR extends VkSubpassDescription2
pub type FragmentShadingRateAttachmentInfoKHR = C.VkFragmentShadingRateAttachmentInfoKHR

@[typedef]
pub struct C.VkFragmentShadingRateAttachmentInfoKHR {
pub mut:
	sType                          StructureType = StructureType.fragment_shading_rate_attachment_info_khr
	pNext                          voidptr       = unsafe { nil }
	pFragmentShadingRateAttachment &AttachmentReference2
	shadingRateAttachmentTexelSize Extent2D
}

// PipelineFragmentShadingRateStateCreateInfoKHR extends VkGraphicsPipelineCreateInfo
pub type PipelineFragmentShadingRateStateCreateInfoKHR = C.VkPipelineFragmentShadingRateStateCreateInfoKHR

@[typedef]
pub struct C.VkPipelineFragmentShadingRateStateCreateInfoKHR {
pub mut:
	sType        StructureType = StructureType.pipeline_fragment_shading_rate_state_create_info_khr
	pNext        voidptr       = unsafe { nil }
	fragmentSize Extent2D
	combinerOps  [2]FragmentShadingRateCombinerOpKHR
}

// PhysicalDeviceFragmentShadingRateFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceFragmentShadingRateFeaturesKHR = C.VkPhysicalDeviceFragmentShadingRateFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceFragmentShadingRateFeaturesKHR {
pub mut:
	sType                         StructureType = StructureType.physical_device_fragment_shading_rate_features_khr
	pNext                         voidptr       = unsafe { nil }
	pipelineFragmentShadingRate   Bool32
	primitiveFragmentShadingRate  Bool32
	attachmentFragmentShadingRate Bool32
}

// PhysicalDeviceFragmentShadingRatePropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceFragmentShadingRatePropertiesKHR = C.VkPhysicalDeviceFragmentShadingRatePropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceFragmentShadingRatePropertiesKHR {
pub mut:
	sType                                                StructureType = StructureType.physical_device_fragment_shading_rate_properties_khr
	pNext                                                voidptr       = unsafe { nil }
	minFragmentShadingRateAttachmentTexelSize            Extent2D
	maxFragmentShadingRateAttachmentTexelSize            Extent2D
	maxFragmentShadingRateAttachmentTexelSizeAspectRatio u32
	primitiveFragmentShadingRateWithMultipleViewports    Bool32
	layeredShadingRateAttachments                        Bool32
	fragmentShadingRateNonTrivialCombinerOps             Bool32
	maxFragmentSize                                      Extent2D
	maxFragmentSizeAspectRatio                           u32
	maxFragmentShadingRateCoverageSamples                u32
	maxFragmentShadingRateRasterizationSamples           SampleCountFlagBits
	fragmentShadingRateWithShaderDepthStencilWrites      Bool32
	fragmentShadingRateWithSampleMask                    Bool32
	fragmentShadingRateWithShaderSampleMask              Bool32
	fragmentShadingRateWithConservativeRasterization     Bool32
	fragmentShadingRateWithFragmentShaderInterlock       Bool32
	fragmentShadingRateWithCustomSampleLocations         Bool32
	fragmentShadingRateStrictMultiplyCombiner            Bool32
}

pub type PhysicalDeviceFragmentShadingRateKHR = C.VkPhysicalDeviceFragmentShadingRateKHR

@[typedef]
pub struct C.VkPhysicalDeviceFragmentShadingRateKHR {
pub mut:
	sType        StructureType = StructureType.physical_device_fragment_shading_rate_khr
	pNext        voidptr       = unsafe { nil }
	sampleCounts SampleCountFlags
	fragmentSize Extent2D
}

// RenderingFragmentShadingRateAttachmentInfoKHR extends VkRenderingInfo
pub type RenderingFragmentShadingRateAttachmentInfoKHR = C.VkRenderingFragmentShadingRateAttachmentInfoKHR

@[typedef]
pub struct C.VkRenderingFragmentShadingRateAttachmentInfoKHR {
pub mut:
	sType                          StructureType = StructureType.rendering_fragment_shading_rate_attachment_info_khr
	pNext                          voidptr       = unsafe { nil }
	imageView                      ImageView
	imageLayout                    ImageLayout
	shadingRateAttachmentTexelSize Extent2D
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceFragmentShadingRatesKHR(physical_device PhysicalDevice, p_fragment_shading_rate_count &u32, mut p_fragment_shading_rates PhysicalDeviceFragmentShadingRateKHR) Result

pub type PFN_vkGetPhysicalDeviceFragmentShadingRatesKHR = fn (physical_device PhysicalDevice, p_fragment_shading_rate_count &u32, mut p_fragment_shading_rates PhysicalDeviceFragmentShadingRateKHR) Result

@[inline]
pub fn get_physical_device_fragment_shading_rates_khr(physical_device PhysicalDevice,
	p_fragment_shading_rate_count &u32,
	mut p_fragment_shading_rates PhysicalDeviceFragmentShadingRateKHR) Result {
	return C.vkGetPhysicalDeviceFragmentShadingRatesKHR(physical_device, p_fragment_shading_rate_count, mut
		p_fragment_shading_rates)
}

/*@[keep_args_alive]
fn C.vkCmdSetFragmentShadingRateKHR(
 command_buffer CommandBuffer,  p_fragment_size &Extent2D,  combiner_ops [2]FragmentShadingRateCombinerOpKHR)
pub type PFN_vkCmdSetFragmentShadingRateKHR = fn(command_buffer CommandBuffer, p_fragment_size &Extent2D, combiner_ops [2]FragmentShadingRateCombinerOpKHR)
@[inline]
pub fn cmd_set_fragment_shading_rate_khr(
command_buffer CommandBuffer,
p_fragment_size &Extent2D,
combiner_ops [2]FragmentShadingRateCombinerOpKHR) {
    C.vkCmdSetFragmentShadingRateKHR( command_buffer, p_fragment_size, combiner_ops)
}

*/

pub const khr_dynamic_rendering_local_read_spec_version = 1
pub const khr_dynamic_rendering_local_read_extension_name = c'VK_KHR_dynamic_rendering_local_read'

pub type PhysicalDeviceDynamicRenderingLocalReadFeaturesKHR = C.VkPhysicalDeviceDynamicRenderingLocalReadFeatures

pub type RenderingAttachmentLocationInfoKHR = C.VkRenderingAttachmentLocationInfo

pub type RenderingInputAttachmentIndexInfoKHR = C.VkRenderingInputAttachmentIndexInfo

@[keep_args_alive]
fn C.vkCmdSetRenderingAttachmentLocationsKHR(command_buffer CommandBuffer, p_location_info &RenderingAttachmentLocationInfo)

pub type PFN_vkCmdSetRenderingAttachmentLocationsKHR = fn (command_buffer CommandBuffer, p_location_info &RenderingAttachmentLocationInfo)

@[inline]
pub fn cmd_set_rendering_attachment_locations_khr(command_buffer CommandBuffer,
	p_location_info &RenderingAttachmentLocationInfo) {
	C.vkCmdSetRenderingAttachmentLocationsKHR(command_buffer, p_location_info)
}

@[keep_args_alive]
fn C.vkCmdSetRenderingInputAttachmentIndicesKHR(command_buffer CommandBuffer, p_input_attachment_index_info &RenderingInputAttachmentIndexInfo)

pub type PFN_vkCmdSetRenderingInputAttachmentIndicesKHR = fn (command_buffer CommandBuffer, p_input_attachment_index_info &RenderingInputAttachmentIndexInfo)

@[inline]
pub fn cmd_set_rendering_input_attachment_indices_khr(command_buffer CommandBuffer,
	p_input_attachment_index_info &RenderingInputAttachmentIndexInfo) {
	C.vkCmdSetRenderingInputAttachmentIndicesKHR(command_buffer, p_input_attachment_index_info)
}

pub const khr_shader_quad_control_spec_version = 1
pub const khr_shader_quad_control_extension_name = c'VK_KHR_shader_quad_control'
// PhysicalDeviceShaderQuadControlFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderQuadControlFeaturesKHR = C.VkPhysicalDeviceShaderQuadControlFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceShaderQuadControlFeaturesKHR {
pub mut:
	sType             StructureType = StructureType.physical_device_shader_quad_control_features_khr
	pNext             voidptr       = unsafe { nil }
	shaderQuadControl Bool32
}

pub const khr_spirv_1_4_spec_version = 1
pub const khr_spirv_1_4_extension_name = c'VK_KHR_spirv_1_4'

pub const khr_surface_protected_capabilities_spec_version = 1
pub const khr_surface_protected_capabilities_extension_name = c'VK_KHR_surface_protected_capabilities'
// SurfaceProtectedCapabilitiesKHR extends VkSurfaceCapabilities2KHR
pub type SurfaceProtectedCapabilitiesKHR = C.VkSurfaceProtectedCapabilitiesKHR

@[typedef]
pub struct C.VkSurfaceProtectedCapabilitiesKHR {
pub mut:
	sType             StructureType = StructureType.surface_protected_capabilities_khr
	pNext             voidptr       = unsafe { nil }
	supportsProtected Bool32
}

pub const khr_separate_depth_stencil_layouts_spec_version = 1
pub const khr_separate_depth_stencil_layouts_extension_name = c'VK_KHR_separate_depth_stencil_layouts'

pub type PhysicalDeviceSeparateDepthStencilLayoutsFeaturesKHR = C.VkPhysicalDeviceSeparateDepthStencilLayoutsFeatures

pub type AttachmentReferenceStencilLayoutKHR = C.VkAttachmentReferenceStencilLayout

pub type AttachmentDescriptionStencilLayoutKHR = C.VkAttachmentDescriptionStencilLayout

pub const khr_present_wait_spec_version = 1
pub const khr_present_wait_extension_name = c'VK_KHR_present_wait'
// PhysicalDevicePresentWaitFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePresentWaitFeaturesKHR = C.VkPhysicalDevicePresentWaitFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDevicePresentWaitFeaturesKHR {
pub mut:
	sType       StructureType = StructureType.physical_device_present_wait_features_khr
	pNext       voidptr       = unsafe { nil }
	presentWait Bool32
}

@[keep_args_alive]
fn C.vkWaitForPresentKHR(device Device, swapchain SwapchainKHR, present_id u64, timeout u64) Result

pub type PFN_vkWaitForPresentKHR = fn (device Device, swapchain SwapchainKHR, present_id u64, timeout u64) Result

@[inline]
pub fn wait_for_present_khr(device Device,
	swapchain SwapchainKHR,
	present_id u64,
	timeout u64) Result {
	return C.vkWaitForPresentKHR(device, swapchain, present_id, timeout)
}

pub const khr_uniform_buffer_standard_layout_spec_version = 1
pub const khr_uniform_buffer_standard_layout_extension_name = c'VK_KHR_uniform_buffer_standard_layout'

pub type PhysicalDeviceUniformBufferStandardLayoutFeaturesKHR = C.VkPhysicalDeviceUniformBufferStandardLayoutFeatures

pub const khr_buffer_device_address_spec_version = 1
pub const khr_buffer_device_address_extension_name = c'VK_KHR_buffer_device_address'

pub type PhysicalDeviceBufferDeviceAddressFeaturesKHR = C.VkPhysicalDeviceBufferDeviceAddressFeatures

pub type BufferDeviceAddressInfoKHR = C.VkBufferDeviceAddressInfo

pub type BufferOpaqueCaptureAddressCreateInfoKHR = C.VkBufferOpaqueCaptureAddressCreateInfo

pub type MemoryOpaqueCaptureAddressAllocateInfoKHR = C.VkMemoryOpaqueCaptureAddressAllocateInfo

pub type DeviceMemoryOpaqueCaptureAddressInfoKHR = C.VkDeviceMemoryOpaqueCaptureAddressInfo

@[keep_args_alive]
fn C.vkGetBufferDeviceAddressKHR(device Device, p_info &BufferDeviceAddressInfo) DeviceAddress

pub type PFN_vkGetBufferDeviceAddressKHR = fn (device Device, p_info &BufferDeviceAddressInfo) DeviceAddress

@[inline]
pub fn get_buffer_device_address_khr(device Device,
	p_info &BufferDeviceAddressInfo) DeviceAddress {
	return C.vkGetBufferDeviceAddressKHR(device, p_info)
}

@[keep_args_alive]
fn C.vkGetBufferOpaqueCaptureAddressKHR(device Device, p_info &BufferDeviceAddressInfo) u64

pub type PFN_vkGetBufferOpaqueCaptureAddressKHR = fn (device Device, p_info &BufferDeviceAddressInfo) u64

@[inline]
pub fn get_buffer_opaque_capture_address_khr(device Device,
	p_info &BufferDeviceAddressInfo) u64 {
	return C.vkGetBufferOpaqueCaptureAddressKHR(device, p_info)
}

@[keep_args_alive]
fn C.vkGetDeviceMemoryOpaqueCaptureAddressKHR(device Device, p_info &DeviceMemoryOpaqueCaptureAddressInfo) u64

pub type PFN_vkGetDeviceMemoryOpaqueCaptureAddressKHR = fn (device Device, p_info &DeviceMemoryOpaqueCaptureAddressInfo) u64

@[inline]
pub fn get_device_memory_opaque_capture_address_khr(device Device,
	p_info &DeviceMemoryOpaqueCaptureAddressInfo) u64 {
	return C.vkGetDeviceMemoryOpaqueCaptureAddressKHR(device, p_info)
}

// Pointer to VkDeferredOperationKHR_T
pub type DeferredOperationKHR = voidptr

pub const khr_deferred_host_operations_spec_version = 4
pub const khr_deferred_host_operations_extension_name = c'VK_KHR_deferred_host_operations'

@[keep_args_alive]
fn C.vkCreateDeferredOperationKHR(device Device, p_allocator &AllocationCallbacks, p_deferred_operation &DeferredOperationKHR) Result

pub type PFN_vkCreateDeferredOperationKHR = fn (device Device, p_allocator &AllocationCallbacks, p_deferred_operation &DeferredOperationKHR) Result

@[inline]
pub fn create_deferred_operation_khr(device Device,
	p_allocator &AllocationCallbacks,
	p_deferred_operation &DeferredOperationKHR) Result {
	return C.vkCreateDeferredOperationKHR(device, p_allocator, p_deferred_operation)
}

@[keep_args_alive]
fn C.vkDestroyDeferredOperationKHR(device Device, operation DeferredOperationKHR, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyDeferredOperationKHR = fn (device Device, operation DeferredOperationKHR, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_deferred_operation_khr(device Device,
	operation DeferredOperationKHR,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyDeferredOperationKHR(device, operation, p_allocator)
}

@[keep_args_alive]
fn C.vkGetDeferredOperationMaxConcurrencyKHR(device Device, operation DeferredOperationKHR) u32

pub type PFN_vkGetDeferredOperationMaxConcurrencyKHR = fn (device Device, operation DeferredOperationKHR) u32

@[inline]
pub fn get_deferred_operation_max_concurrency_khr(device Device,
	operation DeferredOperationKHR) u32 {
	return C.vkGetDeferredOperationMaxConcurrencyKHR(device, operation)
}

@[keep_args_alive]
fn C.vkGetDeferredOperationResultKHR(device Device, operation DeferredOperationKHR) Result

pub type PFN_vkGetDeferredOperationResultKHR = fn (device Device, operation DeferredOperationKHR) Result

@[inline]
pub fn get_deferred_operation_result_khr(device Device,
	operation DeferredOperationKHR) Result {
	return C.vkGetDeferredOperationResultKHR(device, operation)
}

@[keep_args_alive]
fn C.vkDeferredOperationJoinKHR(device Device, operation DeferredOperationKHR) Result

pub type PFN_vkDeferredOperationJoinKHR = fn (device Device, operation DeferredOperationKHR) Result

@[inline]
pub fn deferred_operation_join_khr(device Device,
	operation DeferredOperationKHR) Result {
	return C.vkDeferredOperationJoinKHR(device, operation)
}

pub const khr_pipeline_executable_properties_spec_version = 1
pub const khr_pipeline_executable_properties_extension_name = c'VK_KHR_pipeline_executable_properties'

pub enum PipelineExecutableStatisticFormatKHR as u32 {
	bool32       = 0
	int64        = 1
	uint64       = 2
	float64      = 3
	max_enum_khr = max_int
}
// PhysicalDevicePipelineExecutablePropertiesFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePipelineExecutablePropertiesFeaturesKHR = C.VkPhysicalDevicePipelineExecutablePropertiesFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDevicePipelineExecutablePropertiesFeaturesKHR {
pub mut:
	sType                  StructureType = StructureType.physical_device_pipeline_executable_properties_features_khr
	pNext                  voidptr       = unsafe { nil }
	pipelineExecutableInfo Bool32
}

pub type PipelineInfoKHR = C.VkPipelineInfoKHR

@[typedef]
pub struct C.VkPipelineInfoKHR {
pub mut:
	sType    StructureType = StructureType.pipeline_info_khr
	pNext    voidptr       = unsafe { nil }
	pipeline Pipeline
}

pub type PipelineExecutablePropertiesKHR = C.VkPipelineExecutablePropertiesKHR

@[typedef]
pub struct C.VkPipelineExecutablePropertiesKHR {
pub mut:
	sType        StructureType = StructureType.pipeline_executable_properties_khr
	pNext        voidptr       = unsafe { nil }
	stages       ShaderStageFlags
	name         [max_description_size]char
	description  [max_description_size]char
	subgroupSize u32
}

pub type PipelineExecutableInfoKHR = C.VkPipelineExecutableInfoKHR

@[typedef]
pub struct C.VkPipelineExecutableInfoKHR {
pub mut:
	sType           StructureType = StructureType.pipeline_executable_info_khr
	pNext           voidptr       = unsafe { nil }
	pipeline        Pipeline
	executableIndex u32
}

pub type PipelineExecutableStatisticValueKHR = C.VkPipelineExecutableStatisticValueKHR

@[typedef]
pub union C.VkPipelineExecutableStatisticValueKHR {
pub mut:
	b32 Bool32
	i64 i64
	u64 u64
	f64 f64
}

pub type PipelineExecutableStatisticKHR = C.VkPipelineExecutableStatisticKHR

@[typedef]
pub struct C.VkPipelineExecutableStatisticKHR {
pub mut:
	sType       StructureType = StructureType.pipeline_executable_statistic_khr
	pNext       voidptr       = unsafe { nil }
	name        [max_description_size]char
	description [max_description_size]char
	format      PipelineExecutableStatisticFormatKHR
	value       PipelineExecutableStatisticValueKHR
}

pub type PipelineExecutableInternalRepresentationKHR = C.VkPipelineExecutableInternalRepresentationKHR

@[typedef]
pub struct C.VkPipelineExecutableInternalRepresentationKHR {
pub mut:
	sType       StructureType = StructureType.pipeline_executable_internal_representation_khr
	pNext       voidptr       = unsafe { nil }
	name        [max_description_size]char
	description [max_description_size]char
	isText      Bool32
	dataSize    usize
	pData       voidptr
}

@[keep_args_alive]
fn C.vkGetPipelineExecutablePropertiesKHR(device Device, p_pipeline_info &PipelineInfoKHR, p_executable_count &u32, mut p_properties PipelineExecutablePropertiesKHR) Result

pub type PFN_vkGetPipelineExecutablePropertiesKHR = fn (device Device, p_pipeline_info &PipelineInfoKHR, p_executable_count &u32, mut p_properties PipelineExecutablePropertiesKHR) Result

@[inline]
pub fn get_pipeline_executable_properties_khr(device Device,
	p_pipeline_info &PipelineInfoKHR,
	p_executable_count &u32,
	mut p_properties PipelineExecutablePropertiesKHR) Result {
	return C.vkGetPipelineExecutablePropertiesKHR(device, p_pipeline_info, p_executable_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkGetPipelineExecutableStatisticsKHR(device Device, p_executable_info &PipelineExecutableInfoKHR, p_statistic_count &u32, mut p_statistics PipelineExecutableStatisticKHR) Result

pub type PFN_vkGetPipelineExecutableStatisticsKHR = fn (device Device, p_executable_info &PipelineExecutableInfoKHR, p_statistic_count &u32, mut p_statistics PipelineExecutableStatisticKHR) Result

@[inline]
pub fn get_pipeline_executable_statistics_khr(device Device,
	p_executable_info &PipelineExecutableInfoKHR,
	p_statistic_count &u32,
	mut p_statistics PipelineExecutableStatisticKHR) Result {
	return C.vkGetPipelineExecutableStatisticsKHR(device, p_executable_info, p_statistic_count, mut
		p_statistics)
}

@[keep_args_alive]
fn C.vkGetPipelineExecutableInternalRepresentationsKHR(device Device, p_executable_info &PipelineExecutableInfoKHR, p_internal_representation_count &u32, mut p_internal_representations PipelineExecutableInternalRepresentationKHR) Result

pub type PFN_vkGetPipelineExecutableInternalRepresentationsKHR = fn (device Device, p_executable_info &PipelineExecutableInfoKHR, p_internal_representation_count &u32, mut p_internal_representations PipelineExecutableInternalRepresentationKHR) Result

@[inline]
pub fn get_pipeline_executable_internal_representations_khr(device Device,
	p_executable_info &PipelineExecutableInfoKHR,
	p_internal_representation_count &u32,
	mut p_internal_representations PipelineExecutableInternalRepresentationKHR) Result {
	return C.vkGetPipelineExecutableInternalRepresentationsKHR(device, p_executable_info,
		p_internal_representation_count, mut p_internal_representations)
}

pub const khr_map_memory_2_spec_version = 1
pub const khr_map_memory_2_extension_name = c'VK_KHR_map_memory2'

pub type MemoryUnmapFlagBitsKHR = MemoryUnmapFlagBits

pub type MemoryUnmapFlagsKHR = u32
pub type MemoryMapInfoKHR = C.VkMemoryMapInfo

pub type MemoryUnmapInfoKHR = C.VkMemoryUnmapInfo

@[keep_args_alive]
fn C.vkMapMemory2KHR(device Device, p_memory_map_info &MemoryMapInfo, pp_data &voidptr) Result

pub type PFN_vkMapMemory2KHR = fn (device Device, p_memory_map_info &MemoryMapInfo, pp_data &voidptr) Result

@[inline]
pub fn map_memory2_khr(device Device,
	p_memory_map_info &MemoryMapInfo,
	pp_data &voidptr) Result {
	return C.vkMapMemory2KHR(device, p_memory_map_info, pp_data)
}

@[keep_args_alive]
fn C.vkUnmapMemory2KHR(device Device, p_memory_unmap_info &MemoryUnmapInfo) Result

pub type PFN_vkUnmapMemory2KHR = fn (device Device, p_memory_unmap_info &MemoryUnmapInfo) Result

@[inline]
pub fn unmap_memory2_khr(device Device,
	p_memory_unmap_info &MemoryUnmapInfo) Result {
	return C.vkUnmapMemory2KHR(device, p_memory_unmap_info)
}

pub const khr_shader_integer_dot_product_spec_version = 1
pub const khr_shader_integer_dot_product_extension_name = c'VK_KHR_shader_integer_dot_product'

pub type PhysicalDeviceShaderIntegerDotProductFeaturesKHR = C.VkPhysicalDeviceShaderIntegerDotProductFeatures

pub type PhysicalDeviceShaderIntegerDotProductPropertiesKHR = C.VkPhysicalDeviceShaderIntegerDotProductProperties

pub const khr_pipeline_library_spec_version = 1
pub const khr_pipeline_library_extension_name = c'VK_KHR_pipeline_library'
// PipelineLibraryCreateInfoKHR extends VkGraphicsPipelineCreateInfo
pub type PipelineLibraryCreateInfoKHR = C.VkPipelineLibraryCreateInfoKHR

@[typedef]
pub struct C.VkPipelineLibraryCreateInfoKHR {
pub mut:
	sType        StructureType = StructureType.pipeline_library_create_info_khr
	pNext        voidptr       = unsafe { nil }
	libraryCount u32
	pLibraries   &Pipeline
}

pub const khr_shader_non_semantic_info_spec_version = 1
pub const khr_shader_non_semantic_info_extension_name = c'VK_KHR_shader_non_semantic_info'

pub const khr_present_id_spec_version = 1
pub const khr_present_id_extension_name = c'VK_KHR_present_id'
// PresentIdKHR extends VkPresentInfoKHR
pub type PresentIdKHR = C.VkPresentIdKHR

@[typedef]
pub struct C.VkPresentIdKHR {
pub mut:
	sType          StructureType = StructureType.present_id_khr
	pNext          voidptr       = unsafe { nil }
	swapchainCount u32
	pPresentIds    &u64
}

// PhysicalDevicePresentIdFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePresentIdFeaturesKHR = C.VkPhysicalDevicePresentIdFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDevicePresentIdFeaturesKHR {
pub mut:
	sType     StructureType = StructureType.physical_device_present_id_features_khr
	pNext     voidptr       = unsafe { nil }
	presentId Bool32
}

pub const khr_video_encode_queue_spec_version = 12
pub const khr_video_encode_queue_extension_name = c'VK_KHR_video_encode_queue'

pub enum VideoEncodeTuningModeKHR as u32 {
	default           = 0
	high_quality      = 1
	low_latency       = 2
	ultra_low_latency = 3
	lossless          = 4
	max_enum_khr      = max_int
}

pub enum VideoEncodeFlagBitsKHR as u32 {
	intra_refresh               = u32(0x00000004)
	with_quantization_delta_map = u32(0x00000001)
	with_emphasis_map           = u32(0x00000002)
	max_enum_khr                = max_int
}
pub type VideoEncodeFlagsKHR = u32

pub enum VideoEncodeCapabilityFlagBitsKHR as u32 {
	preceding_externally_encoded_bytes            = u32(0x00000001)
	insufficient_bitstream_buffer_range_detection = u32(0x00000002)
	quantization_delta_map                        = u32(0x00000004)
	emphasis_map                                  = u32(0x00000008)
	max_enum_khr                                  = max_int
}
pub type VideoEncodeCapabilityFlagsKHR = u32

pub enum VideoEncodeRateControlModeFlagBitsKHR as u32 {
	default      = 0
	disabled     = u32(0x00000001)
	cbr          = u32(0x00000002)
	vbr          = u32(0x00000004)
	max_enum_khr = max_int
}
pub type VideoEncodeRateControlModeFlagsKHR = u32

pub enum VideoEncodeFeedbackFlagBitsKHR as u32 {
	bitstream_buffer_offset = u32(0x00000001)
	bitstream_bytes_written = u32(0x00000002)
	bitstream_has_overrides = u32(0x00000004)
	max_enum_khr            = max_int
}
pub type VideoEncodeFeedbackFlagsKHR = u32

pub enum VideoEncodeUsageFlagBitsKHR as u32 {
	default      = 0
	transcoding  = u32(0x00000001)
	streaming    = u32(0x00000002)
	recording    = u32(0x00000004)
	conferencing = u32(0x00000008)
	max_enum_khr = max_int
}
pub type VideoEncodeUsageFlagsKHR = u32

pub enum VideoEncodeContentFlagBitsKHR as u32 {
	default      = 0
	camera       = u32(0x00000001)
	desktop      = u32(0x00000002)
	rendered     = u32(0x00000004)
	max_enum_khr = max_int
}
pub type VideoEncodeContentFlagsKHR = u32
pub type VideoEncodeRateControlFlagsKHR = u32
pub type VideoEncodeInfoKHR = C.VkVideoEncodeInfoKHR

@[typedef]
pub struct C.VkVideoEncodeInfoKHR {
pub mut:
	sType                           StructureType = StructureType.video_encode_info_khr
	pNext                           voidptr       = unsafe { nil }
	flags                           VideoEncodeFlagsKHR
	dstBuffer                       Buffer
	dstBufferOffset                 DeviceSize
	dstBufferRange                  DeviceSize
	srcPictureResource              VideoPictureResourceInfoKHR
	pSetupReferenceSlot             &VideoReferenceSlotInfoKHR
	referenceSlotCount              u32
	pReferenceSlots                 &VideoReferenceSlotInfoKHR
	precedingExternallyEncodedBytes u32
}

// VideoEncodeCapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoEncodeCapabilitiesKHR = C.VkVideoEncodeCapabilitiesKHR

@[typedef]
pub struct C.VkVideoEncodeCapabilitiesKHR {
pub mut:
	sType                         StructureType = StructureType.video_encode_capabilities_khr
	pNext                         voidptr       = unsafe { nil }
	flags                         VideoEncodeCapabilityFlagsKHR
	rateControlModes              VideoEncodeRateControlModeFlagsKHR
	maxRateControlLayers          u32
	maxBitrate                    u64
	maxQualityLevels              u32
	encodeInputPictureGranularity Extent2D
	supportedEncodeFeedbackFlags  VideoEncodeFeedbackFlagsKHR
}

// QueryPoolVideoEncodeFeedbackCreateInfoKHR extends VkQueryPoolCreateInfo
pub type QueryPoolVideoEncodeFeedbackCreateInfoKHR = C.VkQueryPoolVideoEncodeFeedbackCreateInfoKHR

@[typedef]
pub struct C.VkQueryPoolVideoEncodeFeedbackCreateInfoKHR {
pub mut:
	sType               StructureType = StructureType.query_pool_video_encode_feedback_create_info_khr
	pNext               voidptr       = unsafe { nil }
	encodeFeedbackFlags VideoEncodeFeedbackFlagsKHR
}

// VideoEncodeUsageInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub type VideoEncodeUsageInfoKHR = C.VkVideoEncodeUsageInfoKHR

@[typedef]
pub struct C.VkVideoEncodeUsageInfoKHR {
pub mut:
	sType             StructureType = StructureType.video_encode_usage_info_khr
	pNext             voidptr       = unsafe { nil }
	videoUsageHints   VideoEncodeUsageFlagsKHR
	videoContentHints VideoEncodeContentFlagsKHR
	tuningMode        VideoEncodeTuningModeKHR
}

pub type VideoEncodeRateControlLayerInfoKHR = C.VkVideoEncodeRateControlLayerInfoKHR

@[typedef]
pub struct C.VkVideoEncodeRateControlLayerInfoKHR {
pub mut:
	sType                StructureType = StructureType.video_encode_rate_control_layer_info_khr
	pNext                voidptr       = unsafe { nil }
	averageBitrate       u64
	maxBitrate           u64
	frameRateNumerator   u32
	frameRateDenominator u32
}

// VideoEncodeRateControlInfoKHR extends VkVideoCodingControlInfoKHR,VkVideoBeginCodingInfoKHR
pub type VideoEncodeRateControlInfoKHR = C.VkVideoEncodeRateControlInfoKHR

@[typedef]
pub struct C.VkVideoEncodeRateControlInfoKHR {
pub mut:
	sType                        StructureType = StructureType.video_encode_rate_control_info_khr
	pNext                        voidptr       = unsafe { nil }
	flags                        VideoEncodeRateControlFlagsKHR
	rateControlMode              VideoEncodeRateControlModeFlagBitsKHR
	layerCount                   u32
	pLayers                      &VideoEncodeRateControlLayerInfoKHR
	virtualBufferSizeInMs        u32
	initialVirtualBufferSizeInMs u32
}

pub type PhysicalDeviceVideoEncodeQualityLevelInfoKHR = C.VkPhysicalDeviceVideoEncodeQualityLevelInfoKHR

@[typedef]
pub struct C.VkPhysicalDeviceVideoEncodeQualityLevelInfoKHR {
pub mut:
	sType         StructureType = StructureType.physical_device_video_encode_quality_level_info_khr
	pNext         voidptr       = unsafe { nil }
	pVideoProfile &VideoProfileInfoKHR
	qualityLevel  u32
}

pub type VideoEncodeQualityLevelPropertiesKHR = C.VkVideoEncodeQualityLevelPropertiesKHR

@[typedef]
pub struct C.VkVideoEncodeQualityLevelPropertiesKHR {
pub mut:
	sType                          StructureType = StructureType.video_encode_quality_level_properties_khr
	pNext                          voidptr       = unsafe { nil }
	preferredRateControlMode       VideoEncodeRateControlModeFlagBitsKHR
	preferredRateControlLayerCount u32
}

// VideoEncodeQualityLevelInfoKHR extends VkVideoCodingControlInfoKHR,VkVideoSessionParametersCreateInfoKHR
pub type VideoEncodeQualityLevelInfoKHR = C.VkVideoEncodeQualityLevelInfoKHR

@[typedef]
pub struct C.VkVideoEncodeQualityLevelInfoKHR {
pub mut:
	sType        StructureType = StructureType.video_encode_quality_level_info_khr
	pNext        voidptr       = unsafe { nil }
	qualityLevel u32
}

pub type VideoEncodeSessionParametersGetInfoKHR = C.VkVideoEncodeSessionParametersGetInfoKHR

@[typedef]
pub struct C.VkVideoEncodeSessionParametersGetInfoKHR {
pub mut:
	sType                  StructureType = StructureType.video_encode_session_parameters_get_info_khr
	pNext                  voidptr       = unsafe { nil }
	videoSessionParameters VideoSessionParametersKHR
}

pub type VideoEncodeSessionParametersFeedbackInfoKHR = C.VkVideoEncodeSessionParametersFeedbackInfoKHR

@[typedef]
pub struct C.VkVideoEncodeSessionParametersFeedbackInfoKHR {
pub mut:
	sType        StructureType = StructureType.video_encode_session_parameters_feedback_info_khr
	pNext        voidptr       = unsafe { nil }
	hasOverrides Bool32
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceVideoEncodeQualityLevelPropertiesKHR(physical_device PhysicalDevice, p_quality_level_info &PhysicalDeviceVideoEncodeQualityLevelInfoKHR, mut p_quality_level_properties VideoEncodeQualityLevelPropertiesKHR) Result

pub type PFN_vkGetPhysicalDeviceVideoEncodeQualityLevelPropertiesKHR = fn (physical_device PhysicalDevice, p_quality_level_info &PhysicalDeviceVideoEncodeQualityLevelInfoKHR, mut p_quality_level_properties VideoEncodeQualityLevelPropertiesKHR) Result

@[inline]
pub fn get_physical_device_video_encode_quality_level_properties_khr(physical_device PhysicalDevice,
	p_quality_level_info &PhysicalDeviceVideoEncodeQualityLevelInfoKHR,
	mut p_quality_level_properties VideoEncodeQualityLevelPropertiesKHR) Result {
	return C.vkGetPhysicalDeviceVideoEncodeQualityLevelPropertiesKHR(physical_device,
		p_quality_level_info, mut p_quality_level_properties)
}

@[keep_args_alive]
fn C.vkGetEncodedVideoSessionParametersKHR(device Device, p_video_session_parameters_info &VideoEncodeSessionParametersGetInfoKHR, mut p_feedback_info VideoEncodeSessionParametersFeedbackInfoKHR, p_data_size &usize, p_data voidptr) Result

pub type PFN_vkGetEncodedVideoSessionParametersKHR = fn (device Device, p_video_session_parameters_info &VideoEncodeSessionParametersGetInfoKHR, mut p_feedback_info VideoEncodeSessionParametersFeedbackInfoKHR, p_data_size &usize, p_data voidptr) Result

@[inline]
pub fn get_encoded_video_session_parameters_khr(device Device,
	p_video_session_parameters_info &VideoEncodeSessionParametersGetInfoKHR,
	mut p_feedback_info VideoEncodeSessionParametersFeedbackInfoKHR,
	p_data_size &usize,
	p_data voidptr) Result {
	return C.vkGetEncodedVideoSessionParametersKHR(device, p_video_session_parameters_info, mut
		p_feedback_info, p_data_size, p_data)
}

@[keep_args_alive]
fn C.vkCmdEncodeVideoKHR(command_buffer CommandBuffer, p_encode_info &VideoEncodeInfoKHR)

pub type PFN_vkCmdEncodeVideoKHR = fn (command_buffer CommandBuffer, p_encode_info &VideoEncodeInfoKHR)

@[inline]
pub fn cmd_encode_video_khr(command_buffer CommandBuffer,
	p_encode_info &VideoEncodeInfoKHR) {
	C.vkCmdEncodeVideoKHR(command_buffer, p_encode_info)
}

pub const khr_synchronization_2_spec_version = 1
pub const khr_synchronization_2_extension_name = c'VK_KHR_synchronization2'

pub type PipelineStageFlags2KHR = u64
pub type PipelineStageFlagBits2KHR = u64

pub type AccessFlags2KHR = u64
pub type AccessFlagBits2KHR = u64

pub type SubmitFlagBitsKHR = SubmitFlagBits

pub type SubmitFlagsKHR = u32
pub type MemoryBarrier2KHR = C.VkMemoryBarrier2

pub type BufferMemoryBarrier2KHR = C.VkBufferMemoryBarrier2

pub type ImageMemoryBarrier2KHR = C.VkImageMemoryBarrier2

pub type DependencyInfoKHR = C.VkDependencyInfo

pub type SubmitInfo2KHR = C.VkSubmitInfo2

pub type SemaphoreSubmitInfoKHR = C.VkSemaphoreSubmitInfo

pub type CommandBufferSubmitInfoKHR = C.VkCommandBufferSubmitInfo

pub type PhysicalDeviceSynchronization2FeaturesKHR = C.VkPhysicalDeviceSynchronization2Features

@[keep_args_alive]
fn C.vkCmdSetEvent2KHR(command_buffer CommandBuffer, event Event, p_dependency_info &DependencyInfo)

pub type PFN_vkCmdSetEvent2KHR = fn (command_buffer CommandBuffer, event Event, p_dependency_info &DependencyInfo)

@[inline]
pub fn cmd_set_event2_khr(command_buffer CommandBuffer,
	event Event,
	p_dependency_info &DependencyInfo) {
	C.vkCmdSetEvent2KHR(command_buffer, event, p_dependency_info)
}

@[keep_args_alive]
fn C.vkCmdResetEvent2KHR(command_buffer CommandBuffer, event Event, stage_mask PipelineStageFlags2)

pub type PFN_vkCmdResetEvent2KHR = fn (command_buffer CommandBuffer, event Event, stage_mask PipelineStageFlags2)

@[inline]
pub fn cmd_reset_event2_khr(command_buffer CommandBuffer,
	event Event,
	stage_mask PipelineStageFlags2) {
	C.vkCmdResetEvent2KHR(command_buffer, event, stage_mask)
}

@[keep_args_alive]
fn C.vkCmdWaitEvents2KHR(command_buffer CommandBuffer, event_count u32, p_events &Event, p_dependency_infos &DependencyInfo)

pub type PFN_vkCmdWaitEvents2KHR = fn (command_buffer CommandBuffer, event_count u32, p_events &Event, p_dependency_infos &DependencyInfo)

@[inline]
pub fn cmd_wait_events2_khr(command_buffer CommandBuffer,
	event_count u32,
	p_events &Event,
	p_dependency_infos &DependencyInfo) {
	C.vkCmdWaitEvents2KHR(command_buffer, event_count, p_events, p_dependency_infos)
}

@[keep_args_alive]
fn C.vkCmdPipelineBarrier2KHR(command_buffer CommandBuffer, p_dependency_info &DependencyInfo)

pub type PFN_vkCmdPipelineBarrier2KHR = fn (command_buffer CommandBuffer, p_dependency_info &DependencyInfo)

@[inline]
pub fn cmd_pipeline_barrier2_khr(command_buffer CommandBuffer,
	p_dependency_info &DependencyInfo) {
	C.vkCmdPipelineBarrier2KHR(command_buffer, p_dependency_info)
}

@[keep_args_alive]
fn C.vkCmdWriteTimestamp2KHR(command_buffer CommandBuffer, stage PipelineStageFlags2, query_pool QueryPool, query u32)

pub type PFN_vkCmdWriteTimestamp2KHR = fn (command_buffer CommandBuffer, stage PipelineStageFlags2, query_pool QueryPool, query u32)

@[inline]
pub fn cmd_write_timestamp2_khr(command_buffer CommandBuffer,
	stage PipelineStageFlags2,
	query_pool QueryPool,
	query u32) {
	C.vkCmdWriteTimestamp2KHR(command_buffer, stage, query_pool, query)
}

@[keep_args_alive]
fn C.vkQueueSubmit2KHR(queue Queue, submit_count u32, p_submits &SubmitInfo2, fence Fence) Result

pub type PFN_vkQueueSubmit2KHR = fn (queue Queue, submit_count u32, p_submits &SubmitInfo2, fence Fence) Result

@[inline]
pub fn queue_submit2_khr(queue Queue,
	submit_count u32,
	p_submits &SubmitInfo2,
	fence Fence) Result {
	return C.vkQueueSubmit2KHR(queue, submit_count, p_submits, fence)
}

pub const khr_fragment_shader_barycentric_spec_version = 1
pub const khr_fragment_shader_barycentric_extension_name = c'VK_KHR_fragment_shader_barycentric'
// PhysicalDeviceFragmentShaderBarycentricFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceFragmentShaderBarycentricFeaturesKHR = C.VkPhysicalDeviceFragmentShaderBarycentricFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceFragmentShaderBarycentricFeaturesKHR {
pub mut:
	sType                     StructureType = StructureType.physical_device_fragment_shader_barycentric_features_khr
	pNext                     voidptr       = unsafe { nil }
	fragmentShaderBarycentric Bool32
}

// PhysicalDeviceFragmentShaderBarycentricPropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceFragmentShaderBarycentricPropertiesKHR = C.VkPhysicalDeviceFragmentShaderBarycentricPropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceFragmentShaderBarycentricPropertiesKHR {
pub mut:
	sType                                           StructureType = StructureType.physical_device_fragment_shader_barycentric_properties_khr
	pNext                                           voidptr       = unsafe { nil }
	triStripVertexOrderIndependentOfProvokingVertex Bool32
}

pub const khr_shader_subgroup_uniform_control_flow_spec_version = 1
pub const khr_shader_subgroup_uniform_control_flow_extension_name = c'VK_KHR_shader_subgroup_uniform_control_flow'
// PhysicalDeviceShaderSubgroupUniformControlFlowFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderSubgroupUniformControlFlowFeaturesKHR = C.VkPhysicalDeviceShaderSubgroupUniformControlFlowFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceShaderSubgroupUniformControlFlowFeaturesKHR {
pub mut:
	sType                            StructureType = StructureType.physical_device_shader_subgroup_uniform_control_flow_features_khr
	pNext                            voidptr       = unsafe { nil }
	shaderSubgroupUniformControlFlow Bool32
}

pub const khr_zero_initialize_workgroup_memory_spec_version = 1
pub const khr_zero_initialize_workgroup_memory_extension_name = c'VK_KHR_zero_initialize_workgroup_memory'

pub type PhysicalDeviceZeroInitializeWorkgroupMemoryFeaturesKHR = C.VkPhysicalDeviceZeroInitializeWorkgroupMemoryFeatures

pub const khr_workgroup_memory_explicit_layout_spec_version = 1
pub const khr_workgroup_memory_explicit_layout_extension_name = c'VK_KHR_workgroup_memory_explicit_layout'
// PhysicalDeviceWorkgroupMemoryExplicitLayoutFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceWorkgroupMemoryExplicitLayoutFeaturesKHR = C.VkPhysicalDeviceWorkgroupMemoryExplicitLayoutFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceWorkgroupMemoryExplicitLayoutFeaturesKHR {
pub mut:
	sType                                          StructureType = StructureType.physical_device_workgroup_memory_explicit_layout_features_khr
	pNext                                          voidptr       = unsafe { nil }
	workgroupMemoryExplicitLayout                  Bool32
	workgroupMemoryExplicitLayoutScalarBlockLayout Bool32
	workgroupMemoryExplicitLayout8BitAccess        Bool32
	workgroupMemoryExplicitLayout16BitAccess       Bool32
}

pub const khr_copy_commands_2_spec_version = 1
pub const khr_copy_commands_2_extension_name = c'VK_KHR_copy_commands2'

pub type CopyBufferInfo2KHR = C.VkCopyBufferInfo2

pub type CopyImageInfo2KHR = C.VkCopyImageInfo2

pub type CopyBufferToImageInfo2KHR = C.VkCopyBufferToImageInfo2

pub type CopyImageToBufferInfo2KHR = C.VkCopyImageToBufferInfo2

pub type BlitImageInfo2KHR = C.VkBlitImageInfo2

pub type ResolveImageInfo2KHR = C.VkResolveImageInfo2

pub type BufferCopy2KHR = C.VkBufferCopy2

pub type ImageCopy2KHR = C.VkImageCopy2

pub type ImageBlit2KHR = C.VkImageBlit2

pub type BufferImageCopy2KHR = C.VkBufferImageCopy2

pub type ImageResolve2KHR = C.VkImageResolve2

@[keep_args_alive]
fn C.vkCmdCopyBuffer2KHR(command_buffer CommandBuffer, p_copy_buffer_info &CopyBufferInfo2)

pub type PFN_vkCmdCopyBuffer2KHR = fn (command_buffer CommandBuffer, p_copy_buffer_info &CopyBufferInfo2)

@[inline]
pub fn cmd_copy_buffer2_khr(command_buffer CommandBuffer,
	p_copy_buffer_info &CopyBufferInfo2) {
	C.vkCmdCopyBuffer2KHR(command_buffer, p_copy_buffer_info)
}

@[keep_args_alive]
fn C.vkCmdCopyImage2KHR(command_buffer CommandBuffer, p_copy_image_info &CopyImageInfo2)

pub type PFN_vkCmdCopyImage2KHR = fn (command_buffer CommandBuffer, p_copy_image_info &CopyImageInfo2)

@[inline]
pub fn cmd_copy_image2_khr(command_buffer CommandBuffer,
	p_copy_image_info &CopyImageInfo2) {
	C.vkCmdCopyImage2KHR(command_buffer, p_copy_image_info)
}

@[keep_args_alive]
fn C.vkCmdCopyBufferToImage2KHR(command_buffer CommandBuffer, p_copy_buffer_to_image_info &CopyBufferToImageInfo2)

pub type PFN_vkCmdCopyBufferToImage2KHR = fn (command_buffer CommandBuffer, p_copy_buffer_to_image_info &CopyBufferToImageInfo2)

@[inline]
pub fn cmd_copy_buffer_to_image2_khr(command_buffer CommandBuffer,
	p_copy_buffer_to_image_info &CopyBufferToImageInfo2) {
	C.vkCmdCopyBufferToImage2KHR(command_buffer, p_copy_buffer_to_image_info)
}

@[keep_args_alive]
fn C.vkCmdCopyImageToBuffer2KHR(command_buffer CommandBuffer, p_copy_image_to_buffer_info &CopyImageToBufferInfo2)

pub type PFN_vkCmdCopyImageToBuffer2KHR = fn (command_buffer CommandBuffer, p_copy_image_to_buffer_info &CopyImageToBufferInfo2)

@[inline]
pub fn cmd_copy_image_to_buffer2_khr(command_buffer CommandBuffer,
	p_copy_image_to_buffer_info &CopyImageToBufferInfo2) {
	C.vkCmdCopyImageToBuffer2KHR(command_buffer, p_copy_image_to_buffer_info)
}

@[keep_args_alive]
fn C.vkCmdBlitImage2KHR(command_buffer CommandBuffer, p_blit_image_info &BlitImageInfo2)

pub type PFN_vkCmdBlitImage2KHR = fn (command_buffer CommandBuffer, p_blit_image_info &BlitImageInfo2)

@[inline]
pub fn cmd_blit_image2_khr(command_buffer CommandBuffer,
	p_blit_image_info &BlitImageInfo2) {
	C.vkCmdBlitImage2KHR(command_buffer, p_blit_image_info)
}

@[keep_args_alive]
fn C.vkCmdResolveImage2KHR(command_buffer CommandBuffer, p_resolve_image_info &ResolveImageInfo2)

pub type PFN_vkCmdResolveImage2KHR = fn (command_buffer CommandBuffer, p_resolve_image_info &ResolveImageInfo2)

@[inline]
pub fn cmd_resolve_image2_khr(command_buffer CommandBuffer,
	p_resolve_image_info &ResolveImageInfo2) {
	C.vkCmdResolveImage2KHR(command_buffer, p_resolve_image_info)
}

pub const khr_format_feature_flags_2_spec_version = 2
pub const khr_format_feature_flags_2_extension_name = c'VK_KHR_format_feature_flags2'

pub type FormatFeatureFlags2KHR = u64
pub type FormatFeatureFlagBits2KHR = u64

pub type FormatProperties3KHR = C.VkFormatProperties3

pub const khr_ray_tracing_maintenance_1_spec_version = 1
pub const khr_ray_tracing_maintenance_1_extension_name = c'VK_KHR_ray_tracing_maintenance1'
// PhysicalDeviceRayTracingMaintenance1FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRayTracingMaintenance1FeaturesKHR = C.VkPhysicalDeviceRayTracingMaintenance1FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceRayTracingMaintenance1FeaturesKHR {
pub mut:
	sType                                StructureType = StructureType.physical_device_ray_tracing_maintenance1_features_khr
	pNext                                voidptr       = unsafe { nil }
	rayTracingMaintenance1               Bool32
	rayTracingPipelineTraceRaysIndirect2 Bool32
}

pub type TraceRaysIndirectCommand2KHR = C.VkTraceRaysIndirectCommand2KHR

@[typedef]
pub struct C.VkTraceRaysIndirectCommand2KHR {
pub mut:
	raygenShaderRecordAddress         DeviceAddress
	raygenShaderRecordSize            DeviceSize
	missShaderBindingTableAddress     DeviceAddress
	missShaderBindingTableSize        DeviceSize
	missShaderBindingTableStride      DeviceSize
	hitShaderBindingTableAddress      DeviceAddress
	hitShaderBindingTableSize         DeviceSize
	hitShaderBindingTableStride       DeviceSize
	callableShaderBindingTableAddress DeviceAddress
	callableShaderBindingTableSize    DeviceSize
	callableShaderBindingTableStride  DeviceSize
	width                             u32
	height                            u32
	depth                             u32
}

@[keep_args_alive]
fn C.vkCmdTraceRaysIndirect2KHR(command_buffer CommandBuffer, indirect_device_address DeviceAddress)

pub type PFN_vkCmdTraceRaysIndirect2KHR = fn (command_buffer CommandBuffer, indirect_device_address DeviceAddress)

@[inline]
pub fn cmd_trace_rays_indirect2_khr(command_buffer CommandBuffer,
	indirect_device_address DeviceAddress) {
	C.vkCmdTraceRaysIndirect2KHR(command_buffer, indirect_device_address)
}

pub const khr_shader_untyped_pointers_spec_version = 1
pub const khr_shader_untyped_pointers_extension_name = c'VK_KHR_shader_untyped_pointers'
// PhysicalDeviceShaderUntypedPointersFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderUntypedPointersFeaturesKHR = C.VkPhysicalDeviceShaderUntypedPointersFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceShaderUntypedPointersFeaturesKHR {
pub mut:
	sType                 StructureType = StructureType.physical_device_shader_untyped_pointers_features_khr
	pNext                 voidptr       = unsafe { nil }
	shaderUntypedPointers Bool32
}

pub const khr_portability_enumeration_spec_version = 1
pub const khr_portability_enumeration_extension_name = c'VK_KHR_portability_enumeration'

pub const khr_maintenance_4_spec_version = 2
pub const khr_maintenance_4_extension_name = c'VK_KHR_maintenance4'

pub type PhysicalDeviceMaintenance4FeaturesKHR = C.VkPhysicalDeviceMaintenance4Features

pub type PhysicalDeviceMaintenance4PropertiesKHR = C.VkPhysicalDeviceMaintenance4Properties

pub type DeviceBufferMemoryRequirementsKHR = C.VkDeviceBufferMemoryRequirements

pub type DeviceImageMemoryRequirementsKHR = C.VkDeviceImageMemoryRequirements

@[keep_args_alive]
fn C.vkGetDeviceBufferMemoryRequirementsKHR(device Device, p_info &DeviceBufferMemoryRequirements, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetDeviceBufferMemoryRequirementsKHR = fn (device Device, p_info &DeviceBufferMemoryRequirements, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_device_buffer_memory_requirements_khr(device Device,
	p_info &DeviceBufferMemoryRequirements,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetDeviceBufferMemoryRequirementsKHR(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetDeviceImageMemoryRequirementsKHR(device Device, p_info &DeviceImageMemoryRequirements, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetDeviceImageMemoryRequirementsKHR = fn (device Device, p_info &DeviceImageMemoryRequirements, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_device_image_memory_requirements_khr(device Device,
	p_info &DeviceImageMemoryRequirements,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetDeviceImageMemoryRequirementsKHR(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkGetDeviceImageSparseMemoryRequirementsKHR(device Device, p_info &DeviceImageMemoryRequirements, p_sparse_memory_requirement_count &u32, mut p_sparse_memory_requirements SparseImageMemoryRequirements2)

pub type PFN_vkGetDeviceImageSparseMemoryRequirementsKHR = fn (device Device, p_info &DeviceImageMemoryRequirements, p_sparse_memory_requirement_count &u32, mut p_sparse_memory_requirements SparseImageMemoryRequirements2)

@[inline]
pub fn get_device_image_sparse_memory_requirements_khr(device Device,
	p_info &DeviceImageMemoryRequirements,
	p_sparse_memory_requirement_count &u32,
	mut p_sparse_memory_requirements SparseImageMemoryRequirements2) {
	C.vkGetDeviceImageSparseMemoryRequirementsKHR(device, p_info, p_sparse_memory_requirement_count, mut
		p_sparse_memory_requirements)
}

pub const khr_shader_subgroup_rotate_spec_version = 2
pub const khr_shader_subgroup_rotate_extension_name = c'VK_KHR_shader_subgroup_rotate'

pub type PhysicalDeviceShaderSubgroupRotateFeaturesKHR = C.VkPhysicalDeviceShaderSubgroupRotateFeatures

pub const khr_shader_maximal_reconvergence_spec_version = 1
pub const khr_shader_maximal_reconvergence_extension_name = c'VK_KHR_shader_maximal_reconvergence'
// PhysicalDeviceShaderMaximalReconvergenceFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderMaximalReconvergenceFeaturesKHR = C.VkPhysicalDeviceShaderMaximalReconvergenceFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceShaderMaximalReconvergenceFeaturesKHR {
pub mut:
	sType                      StructureType = StructureType.physical_device_shader_maximal_reconvergence_features_khr
	pNext                      voidptr       = unsafe { nil }
	shaderMaximalReconvergence Bool32
}

pub const khr_maintenance_5_spec_version = 1
pub const khr_maintenance_5_extension_name = c'VK_KHR_maintenance5'

pub type PipelineCreateFlags2KHR = u64
pub type PipelineCreateFlagBits2KHR = u64

pub type BufferUsageFlags2KHR = u64
pub type BufferUsageFlagBits2KHR = u64

pub type PhysicalDeviceMaintenance5FeaturesKHR = C.VkPhysicalDeviceMaintenance5Features

pub type PhysicalDeviceMaintenance5PropertiesKHR = C.VkPhysicalDeviceMaintenance5Properties

pub type RenderingAreaInfoKHR = C.VkRenderingAreaInfo

pub type DeviceImageSubresourceInfoKHR = C.VkDeviceImageSubresourceInfo

pub type ImageSubresource2KHR = C.VkImageSubresource2

pub type SubresourceLayout2KHR = C.VkSubresourceLayout2

pub type PipelineCreateFlags2CreateInfoKHR = C.VkPipelineCreateFlags2CreateInfo

pub type BufferUsageFlags2CreateInfoKHR = C.VkBufferUsageFlags2CreateInfo

@[keep_args_alive]
fn C.vkCmdBindIndexBuffer2KHR(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, size DeviceSize, index_type IndexType)

pub type PFN_vkCmdBindIndexBuffer2KHR = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, size DeviceSize, index_type IndexType)

@[inline]
pub fn cmd_bind_index_buffer2_khr(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	size DeviceSize,
	index_type IndexType) {
	C.vkCmdBindIndexBuffer2KHR(command_buffer, buffer, offset, size, index_type)
}

@[keep_args_alive]
fn C.vkGetRenderingAreaGranularityKHR(device Device, p_rendering_area_info &RenderingAreaInfo, mut p_granularity Extent2D)

pub type PFN_vkGetRenderingAreaGranularityKHR = fn (device Device, p_rendering_area_info &RenderingAreaInfo, mut p_granularity Extent2D)

@[inline]
pub fn get_rendering_area_granularity_khr(device Device,
	p_rendering_area_info &RenderingAreaInfo,
	mut p_granularity Extent2D) {
	C.vkGetRenderingAreaGranularityKHR(device, p_rendering_area_info, mut p_granularity)
}

@[keep_args_alive]
fn C.vkGetDeviceImageSubresourceLayoutKHR(device Device, p_info &DeviceImageSubresourceInfo, mut p_layout SubresourceLayout2)

pub type PFN_vkGetDeviceImageSubresourceLayoutKHR = fn (device Device, p_info &DeviceImageSubresourceInfo, mut p_layout SubresourceLayout2)

@[inline]
pub fn get_device_image_subresource_layout_khr(device Device,
	p_info &DeviceImageSubresourceInfo,
	mut p_layout SubresourceLayout2) {
	C.vkGetDeviceImageSubresourceLayoutKHR(device, p_info, mut p_layout)
}

@[keep_args_alive]
fn C.vkGetImageSubresourceLayout2KHR(device Device, image Image, p_subresource &ImageSubresource2, mut p_layout SubresourceLayout2)

pub type PFN_vkGetImageSubresourceLayout2KHR = fn (device Device, image Image, p_subresource &ImageSubresource2, mut p_layout SubresourceLayout2)

@[inline]
pub fn get_image_subresource_layout2_khr(device Device,
	image Image,
	p_subresource &ImageSubresource2,
	mut p_layout SubresourceLayout2) {
	C.vkGetImageSubresourceLayout2KHR(device, image, p_subresource, mut p_layout)
}

pub const khr_present_id_2_spec_version = 1
pub const khr_present_id_2_extension_name = c'VK_KHR_present_id2'
// SurfaceCapabilitiesPresentId2KHR extends VkSurfaceCapabilities2KHR
pub type SurfaceCapabilitiesPresentId2KHR = C.VkSurfaceCapabilitiesPresentId2KHR

@[typedef]
pub struct C.VkSurfaceCapabilitiesPresentId2KHR {
pub mut:
	sType               StructureType = StructureType.surface_capabilities_present_id2_khr
	pNext               voidptr       = unsafe { nil }
	presentId2Supported Bool32
}

// PresentId2KHR extends VkPresentInfoKHR
pub type PresentId2KHR = C.VkPresentId2KHR

@[typedef]
pub struct C.VkPresentId2KHR {
pub mut:
	sType          StructureType = StructureType.present_id2_khr
	pNext          voidptr       = unsafe { nil }
	swapchainCount u32
	pPresentIds    &u64
}

// PhysicalDevicePresentId2FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePresentId2FeaturesKHR = C.VkPhysicalDevicePresentId2FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDevicePresentId2FeaturesKHR {
pub mut:
	sType      StructureType = StructureType.physical_device_present_id2_features_khr
	pNext      voidptr       = unsafe { nil }
	presentId2 Bool32
}

pub const khr_present_wait_2_spec_version = 1
pub const khr_present_wait_2_extension_name = c'VK_KHR_present_wait2'
// SurfaceCapabilitiesPresentWait2KHR extends VkSurfaceCapabilities2KHR
pub type SurfaceCapabilitiesPresentWait2KHR = C.VkSurfaceCapabilitiesPresentWait2KHR

@[typedef]
pub struct C.VkSurfaceCapabilitiesPresentWait2KHR {
pub mut:
	sType                 StructureType = StructureType.surface_capabilities_present_wait2_khr
	pNext                 voidptr       = unsafe { nil }
	presentWait2Supported Bool32
}

// PhysicalDevicePresentWait2FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePresentWait2FeaturesKHR = C.VkPhysicalDevicePresentWait2FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDevicePresentWait2FeaturesKHR {
pub mut:
	sType        StructureType = StructureType.physical_device_present_wait2_features_khr
	pNext        voidptr       = unsafe { nil }
	presentWait2 Bool32
}

pub type PresentWait2InfoKHR = C.VkPresentWait2InfoKHR

@[typedef]
pub struct C.VkPresentWait2InfoKHR {
pub mut:
	sType     StructureType = StructureType.present_wait2_info_khr
	pNext     voidptr       = unsafe { nil }
	presentId u64
	timeout   u64
}

@[keep_args_alive]
fn C.vkWaitForPresent2KHR(device Device, swapchain SwapchainKHR, p_present_wait2_info &PresentWait2InfoKHR) Result

pub type PFN_vkWaitForPresent2KHR = fn (device Device, swapchain SwapchainKHR, p_present_wait2_info &PresentWait2InfoKHR) Result

@[inline]
pub fn wait_for_present2_khr(device Device,
	swapchain SwapchainKHR,
	p_present_wait2_info &PresentWait2InfoKHR) Result {
	return C.vkWaitForPresent2KHR(device, swapchain, p_present_wait2_info)
}

pub const khr_ray_tracing_position_fetch_spec_version = 1
pub const khr_ray_tracing_position_fetch_extension_name = c'VK_KHR_ray_tracing_position_fetch'
// PhysicalDeviceRayTracingPositionFetchFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRayTracingPositionFetchFeaturesKHR = C.VkPhysicalDeviceRayTracingPositionFetchFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceRayTracingPositionFetchFeaturesKHR {
pub mut:
	sType                   StructureType = StructureType.physical_device_ray_tracing_position_fetch_features_khr
	pNext                   voidptr       = unsafe { nil }
	rayTracingPositionFetch Bool32
}

// Pointer to VkPipelineBinaryKHR_T
pub type PipelineBinaryKHR = voidptr

pub const max_pipeline_binary_key_size_khr = u32(32)
pub const khr_pipeline_binary_spec_version = 1
pub const khr_pipeline_binary_extension_name = c'VK_KHR_pipeline_binary'
// PhysicalDevicePipelineBinaryFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePipelineBinaryFeaturesKHR = C.VkPhysicalDevicePipelineBinaryFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDevicePipelineBinaryFeaturesKHR {
pub mut:
	sType            StructureType = StructureType.physical_device_pipeline_binary_features_khr
	pNext            voidptr       = unsafe { nil }
	pipelineBinaries Bool32
}

// PhysicalDevicePipelineBinaryPropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDevicePipelineBinaryPropertiesKHR = C.VkPhysicalDevicePipelineBinaryPropertiesKHR

@[typedef]
pub struct C.VkPhysicalDevicePipelineBinaryPropertiesKHR {
pub mut:
	sType                                  StructureType = StructureType.physical_device_pipeline_binary_properties_khr
	pNext                                  voidptr       = unsafe { nil }
	pipelineBinaryInternalCache            Bool32
	pipelineBinaryInternalCacheControl     Bool32
	pipelineBinaryPrefersInternalCache     Bool32
	pipelineBinaryPrecompiledInternalCache Bool32
	pipelineBinaryCompressedData           Bool32
}

// DevicePipelineBinaryInternalCacheControlKHR extends VkDeviceCreateInfo
pub type DevicePipelineBinaryInternalCacheControlKHR = C.VkDevicePipelineBinaryInternalCacheControlKHR

@[typedef]
pub struct C.VkDevicePipelineBinaryInternalCacheControlKHR {
pub mut:
	sType                StructureType = StructureType.device_pipeline_binary_internal_cache_control_khr
	pNext                voidptr       = unsafe { nil }
	disableInternalCache Bool32
}

pub type PipelineBinaryKeyKHR = C.VkPipelineBinaryKeyKHR

@[typedef]
pub struct C.VkPipelineBinaryKeyKHR {
pub mut:
	sType   StructureType = StructureType.pipeline_binary_key_khr
	pNext   voidptr       = unsafe { nil }
	keySize u32
	key     [max_pipeline_binary_key_size_khr]u8
}

pub type PipelineBinaryDataKHR = C.VkPipelineBinaryDataKHR

@[typedef]
pub struct C.VkPipelineBinaryDataKHR {
pub mut:
	dataSize usize
	pData    voidptr
}

pub type PipelineBinaryKeysAndDataKHR = C.VkPipelineBinaryKeysAndDataKHR

@[typedef]
pub struct C.VkPipelineBinaryKeysAndDataKHR {
pub mut:
	binaryCount         u32
	pPipelineBinaryKeys &PipelineBinaryKeyKHR
	pPipelineBinaryData &PipelineBinaryDataKHR
}

pub type PipelineCreateInfoKHR = C.VkPipelineCreateInfoKHR

@[typedef]
pub struct C.VkPipelineCreateInfoKHR {
pub mut:
	sType StructureType = StructureType.pipeline_create_info_khr
	pNext voidptr       = unsafe { nil }
}

pub type PipelineBinaryCreateInfoKHR = C.VkPipelineBinaryCreateInfoKHR

@[typedef]
pub struct C.VkPipelineBinaryCreateInfoKHR {
pub mut:
	sType               StructureType = StructureType.pipeline_binary_create_info_khr
	pNext               voidptr       = unsafe { nil }
	pKeysAndDataInfo    &PipelineBinaryKeysAndDataKHR
	pipeline            Pipeline
	pPipelineCreateInfo &PipelineCreateInfoKHR
}

// PipelineBinaryInfoKHR extends VkGraphicsPipelineCreateInfo,VkComputePipelineCreateInfo,VkRayTracingPipelineCreateInfoKHR
pub type PipelineBinaryInfoKHR = C.VkPipelineBinaryInfoKHR

@[typedef]
pub struct C.VkPipelineBinaryInfoKHR {
pub mut:
	sType             StructureType = StructureType.pipeline_binary_info_khr
	pNext             voidptr       = unsafe { nil }
	binaryCount       u32
	pPipelineBinaries &PipelineBinaryKHR
}

pub type ReleaseCapturedPipelineDataInfoKHR = C.VkReleaseCapturedPipelineDataInfoKHR

@[typedef]
pub struct C.VkReleaseCapturedPipelineDataInfoKHR {
pub mut:
	sType    StructureType = StructureType.release_captured_pipeline_data_info_khr
	pNext    voidptr       = unsafe { nil }
	pipeline Pipeline
}

pub type PipelineBinaryDataInfoKHR = C.VkPipelineBinaryDataInfoKHR

@[typedef]
pub struct C.VkPipelineBinaryDataInfoKHR {
pub mut:
	sType          StructureType = StructureType.pipeline_binary_data_info_khr
	pNext          voidptr       = unsafe { nil }
	pipelineBinary PipelineBinaryKHR
}

pub type PipelineBinaryHandlesInfoKHR = C.VkPipelineBinaryHandlesInfoKHR

@[typedef]
pub struct C.VkPipelineBinaryHandlesInfoKHR {
pub mut:
	sType               StructureType = StructureType.pipeline_binary_handles_info_khr
	pNext               voidptr       = unsafe { nil }
	pipelineBinaryCount u32
	pPipelineBinaries   &PipelineBinaryKHR
}

@[keep_args_alive]
fn C.vkCreatePipelineBinariesKHR(device Device, p_create_info &PipelineBinaryCreateInfoKHR, p_allocator &AllocationCallbacks, mut p_binaries PipelineBinaryHandlesInfoKHR) Result

pub type PFN_vkCreatePipelineBinariesKHR = fn (device Device, p_create_info &PipelineBinaryCreateInfoKHR, p_allocator &AllocationCallbacks, mut p_binaries PipelineBinaryHandlesInfoKHR) Result

@[inline]
pub fn create_pipeline_binaries_khr(device Device,
	p_create_info &PipelineBinaryCreateInfoKHR,
	p_allocator &AllocationCallbacks,
	mut p_binaries PipelineBinaryHandlesInfoKHR) Result {
	return C.vkCreatePipelineBinariesKHR(device, p_create_info, p_allocator, mut p_binaries)
}

@[keep_args_alive]
fn C.vkDestroyPipelineBinaryKHR(device Device, pipeline_binary PipelineBinaryKHR, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyPipelineBinaryKHR = fn (device Device, pipeline_binary PipelineBinaryKHR, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_pipeline_binary_khr(device Device,
	pipeline_binary PipelineBinaryKHR,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyPipelineBinaryKHR(device, pipeline_binary, p_allocator)
}

@[keep_args_alive]
fn C.vkGetPipelineKeyKHR(device Device, p_pipeline_create_info &PipelineCreateInfoKHR, mut p_pipeline_key PipelineBinaryKeyKHR) Result

pub type PFN_vkGetPipelineKeyKHR = fn (device Device, p_pipeline_create_info &PipelineCreateInfoKHR, mut p_pipeline_key PipelineBinaryKeyKHR) Result

@[inline]
pub fn get_pipeline_key_khr(device Device,
	p_pipeline_create_info &PipelineCreateInfoKHR,
	mut p_pipeline_key PipelineBinaryKeyKHR) Result {
	return C.vkGetPipelineKeyKHR(device, p_pipeline_create_info, mut p_pipeline_key)
}

@[keep_args_alive]
fn C.vkGetPipelineBinaryDataKHR(device Device, p_info &PipelineBinaryDataInfoKHR, mut p_pipeline_binary_key PipelineBinaryKeyKHR, p_pipeline_binary_data_size &usize, p_pipeline_binary_data voidptr) Result

pub type PFN_vkGetPipelineBinaryDataKHR = fn (device Device, p_info &PipelineBinaryDataInfoKHR, mut p_pipeline_binary_key PipelineBinaryKeyKHR, p_pipeline_binary_data_size &usize, p_pipeline_binary_data voidptr) Result

@[inline]
pub fn get_pipeline_binary_data_khr(device Device,
	p_info &PipelineBinaryDataInfoKHR,
	mut p_pipeline_binary_key PipelineBinaryKeyKHR,
	p_pipeline_binary_data_size &usize,
	p_pipeline_binary_data voidptr) Result {
	return C.vkGetPipelineBinaryDataKHR(device, p_info, mut p_pipeline_binary_key, p_pipeline_binary_data_size,
		p_pipeline_binary_data)
}

@[keep_args_alive]
fn C.vkReleaseCapturedPipelineDataKHR(device Device, p_info &ReleaseCapturedPipelineDataInfoKHR, p_allocator &AllocationCallbacks) Result

pub type PFN_vkReleaseCapturedPipelineDataKHR = fn (device Device, p_info &ReleaseCapturedPipelineDataInfoKHR, p_allocator &AllocationCallbacks) Result

@[inline]
pub fn release_captured_pipeline_data_khr(device Device,
	p_info &ReleaseCapturedPipelineDataInfoKHR,
	p_allocator &AllocationCallbacks) Result {
	return C.vkReleaseCapturedPipelineDataKHR(device, p_info, p_allocator)
}

pub const khr_surface_maintenance_1_spec_version = 1
pub const khr_surface_maintenance_1_extension_name = c'VK_KHR_surface_maintenance1'

pub enum PresentScalingFlagBitsKHR as u32 {
	one_to_one           = u32(0x00000001)
	aspect_ratio_stretch = u32(0x00000002)
	stretch              = u32(0x00000004)
	max_enum_khr         = max_int
}
pub type PresentScalingFlagsKHR = u32

pub enum PresentGravityFlagBitsKHR as u32 {
	min          = u32(0x00000001)
	max          = u32(0x00000002)
	centered     = u32(0x00000004)
	max_enum_khr = max_int
}
pub type PresentGravityFlagsKHR = u32

// SurfacePresentModeKHR extends VkPhysicalDeviceSurfaceInfo2KHR
pub type SurfacePresentModeKHR = C.VkSurfacePresentModeKHR

@[typedef]
pub struct C.VkSurfacePresentModeKHR {
pub mut:
	sType       StructureType = StructureType.surface_present_mode_khr
	pNext       voidptr       = unsafe { nil }
	presentMode PresentModeKHR
}

// SurfacePresentScalingCapabilitiesKHR extends VkSurfaceCapabilities2KHR
pub type SurfacePresentScalingCapabilitiesKHR = C.VkSurfacePresentScalingCapabilitiesKHR

@[typedef]
pub struct C.VkSurfacePresentScalingCapabilitiesKHR {
pub mut:
	sType                    StructureType = StructureType.surface_present_scaling_capabilities_khr
	pNext                    voidptr       = unsafe { nil }
	supportedPresentScaling  PresentScalingFlagsKHR
	supportedPresentGravityX PresentGravityFlagsKHR
	supportedPresentGravityY PresentGravityFlagsKHR
	minScaledImageExtent     Extent2D
	maxScaledImageExtent     Extent2D
}

// SurfacePresentModeCompatibilityKHR extends VkSurfaceCapabilities2KHR
pub type SurfacePresentModeCompatibilityKHR = C.VkSurfacePresentModeCompatibilityKHR

@[typedef]
pub struct C.VkSurfacePresentModeCompatibilityKHR {
pub mut:
	sType            StructureType = StructureType.surface_present_mode_compatibility_khr
	pNext            voidptr       = unsafe { nil }
	presentModeCount u32
	pPresentModes    &PresentModeKHR
}

pub const khr_swapchain_maintenance_1_spec_version = 1
pub const khr_swapchain_maintenance_1_extension_name = c'VK_KHR_swapchain_maintenance1'
// PhysicalDeviceSwapchainMaintenance1FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceSwapchainMaintenance1FeaturesKHR = C.VkPhysicalDeviceSwapchainMaintenance1FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceSwapchainMaintenance1FeaturesKHR {
pub mut:
	sType                 StructureType = StructureType.physical_device_swapchain_maintenance1_features_khr
	pNext                 voidptr       = unsafe { nil }
	swapchainMaintenance1 Bool32
}

// SwapchainPresentFenceInfoKHR extends VkPresentInfoKHR
pub type SwapchainPresentFenceInfoKHR = C.VkSwapchainPresentFenceInfoKHR

@[typedef]
pub struct C.VkSwapchainPresentFenceInfoKHR {
pub mut:
	sType          StructureType = StructureType.swapchain_present_fence_info_khr
	pNext          voidptr       = unsafe { nil }
	swapchainCount u32
	pFences        &Fence
}

// SwapchainPresentModesCreateInfoKHR extends VkSwapchainCreateInfoKHR
pub type SwapchainPresentModesCreateInfoKHR = C.VkSwapchainPresentModesCreateInfoKHR

@[typedef]
pub struct C.VkSwapchainPresentModesCreateInfoKHR {
pub mut:
	sType            StructureType = StructureType.swapchain_present_modes_create_info_khr
	pNext            voidptr       = unsafe { nil }
	presentModeCount u32
	pPresentModes    &PresentModeKHR
}

// SwapchainPresentModeInfoKHR extends VkPresentInfoKHR
pub type SwapchainPresentModeInfoKHR = C.VkSwapchainPresentModeInfoKHR

@[typedef]
pub struct C.VkSwapchainPresentModeInfoKHR {
pub mut:
	sType          StructureType = StructureType.swapchain_present_mode_info_khr
	pNext          voidptr       = unsafe { nil }
	swapchainCount u32
	pPresentModes  &PresentModeKHR
}

// SwapchainPresentScalingCreateInfoKHR extends VkSwapchainCreateInfoKHR
pub type SwapchainPresentScalingCreateInfoKHR = C.VkSwapchainPresentScalingCreateInfoKHR

@[typedef]
pub struct C.VkSwapchainPresentScalingCreateInfoKHR {
pub mut:
	sType           StructureType = StructureType.swapchain_present_scaling_create_info_khr
	pNext           voidptr       = unsafe { nil }
	scalingBehavior PresentScalingFlagsKHR
	presentGravityX PresentGravityFlagsKHR
	presentGravityY PresentGravityFlagsKHR
}

pub type ReleaseSwapchainImagesInfoKHR = C.VkReleaseSwapchainImagesInfoKHR

@[typedef]
pub struct C.VkReleaseSwapchainImagesInfoKHR {
pub mut:
	sType           StructureType = StructureType.release_swapchain_images_info_khr
	pNext           voidptr       = unsafe { nil }
	swapchain       SwapchainKHR
	imageIndexCount u32
	pImageIndices   &u32
}

@[keep_args_alive]
fn C.vkReleaseSwapchainImagesKHR(device Device, p_release_info &ReleaseSwapchainImagesInfoKHR) Result

pub type PFN_vkReleaseSwapchainImagesKHR = fn (device Device, p_release_info &ReleaseSwapchainImagesInfoKHR) Result

@[inline]
pub fn release_swapchain_images_khr(device Device,
	p_release_info &ReleaseSwapchainImagesInfoKHR) Result {
	return C.vkReleaseSwapchainImagesKHR(device, p_release_info)
}

pub const khr_cooperative_matrix_spec_version = 2
pub const khr_cooperative_matrix_extension_name = c'VK_KHR_cooperative_matrix'

pub enum ComponentTypeKHR as u32 {
	float16         = 0
	float32         = 1
	float64         = 2
	sint8           = 3
	sint16          = 4
	sint32          = 5
	sint64          = 6
	uint8           = 7
	uint16          = 8
	uint32          = 9
	uint64          = 10
	bfloat16        = 1000141000
	sint8_packed_nv = 1000491000
	uint8_packed_nv = 1000491001
	float8_e4m3_ext = 1000491002
	float8_e5m2_ext = 1000491003
	max_enum_khr    = max_int
}

pub enum ScopeKHR as u32 {
	device       = 1
	workgroup    = 2
	subgroup     = 3
	queue_family = 5
	max_enum_khr = max_int
}
pub type CooperativeMatrixPropertiesKHR = C.VkCooperativeMatrixPropertiesKHR

@[typedef]
pub struct C.VkCooperativeMatrixPropertiesKHR {
pub mut:
	sType                  StructureType = StructureType.cooperative_matrix_properties_khr
	pNext                  voidptr       = unsafe { nil }
	MSize                  u32
	NSize                  u32
	KSize                  u32
	AType                  ComponentTypeKHR
	BType                  ComponentTypeKHR
	CType                  ComponentTypeKHR
	ResultType             ComponentTypeKHR
	saturatingAccumulation Bool32
	scope                  ScopeKHR
}

// PhysicalDeviceCooperativeMatrixFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCooperativeMatrixFeaturesKHR = C.VkPhysicalDeviceCooperativeMatrixFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceCooperativeMatrixFeaturesKHR {
pub mut:
	sType                               StructureType = StructureType.physical_device_cooperative_matrix_features_khr
	pNext                               voidptr       = unsafe { nil }
	cooperativeMatrix                   Bool32
	cooperativeMatrixRobustBufferAccess Bool32
}

// PhysicalDeviceCooperativeMatrixPropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceCooperativeMatrixPropertiesKHR = C.VkPhysicalDeviceCooperativeMatrixPropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceCooperativeMatrixPropertiesKHR {
pub mut:
	sType                            StructureType = StructureType.physical_device_cooperative_matrix_properties_khr
	pNext                            voidptr       = unsafe { nil }
	cooperativeMatrixSupportedStages ShaderStageFlags
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceCooperativeMatrixPropertiesKHR(physical_device PhysicalDevice, p_property_count &u32, mut p_properties CooperativeMatrixPropertiesKHR) Result

pub type PFN_vkGetPhysicalDeviceCooperativeMatrixPropertiesKHR = fn (physical_device PhysicalDevice, p_property_count &u32, mut p_properties CooperativeMatrixPropertiesKHR) Result

@[inline]
pub fn get_physical_device_cooperative_matrix_properties_khr(physical_device PhysicalDevice,
	p_property_count &u32,
	mut p_properties CooperativeMatrixPropertiesKHR) Result {
	return C.vkGetPhysicalDeviceCooperativeMatrixPropertiesKHR(physical_device, p_property_count, mut
		p_properties)
}

pub const khr_compute_shader_derivatives_spec_version = 1
pub const khr_compute_shader_derivatives_extension_name = c'VK_KHR_compute_shader_derivatives'
// PhysicalDeviceComputeShaderDerivativesFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceComputeShaderDerivativesFeaturesKHR = C.VkPhysicalDeviceComputeShaderDerivativesFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceComputeShaderDerivativesFeaturesKHR {
pub mut:
	sType                        StructureType = StructureType.physical_device_compute_shader_derivatives_features_khr
	pNext                        voidptr       = unsafe { nil }
	computeDerivativeGroupQuads  Bool32
	computeDerivativeGroupLinear Bool32
}

// PhysicalDeviceComputeShaderDerivativesPropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceComputeShaderDerivativesPropertiesKHR = C.VkPhysicalDeviceComputeShaderDerivativesPropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceComputeShaderDerivativesPropertiesKHR {
pub mut:
	sType                        StructureType = StructureType.physical_device_compute_shader_derivatives_properties_khr
	pNext                        voidptr       = unsafe { nil }
	meshAndTaskShaderDerivatives Bool32
}

pub const max_video_av1_references_per_frame_khr = u32(7)
pub const khr_video_decode_av1_spec_version = 1
pub const khr_video_decode_av1_extension_name = c'VK_KHR_video_decode_av1'
// VideoDecodeAV1ProfileInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub type VideoDecodeAV1ProfileInfoKHR = C.VkVideoDecodeAV1ProfileInfoKHR

@[typedef]
pub struct C.VkVideoDecodeAV1ProfileInfoKHR {
pub mut:
	sType            StructureType = StructureType.video_decode_av1_profile_info_khr
	pNext            voidptr       = unsafe { nil }
	stdProfile       StdVideoAV1Profile
	filmGrainSupport Bool32
}

// VideoDecodeAV1CapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoDecodeAV1CapabilitiesKHR = C.VkVideoDecodeAV1CapabilitiesKHR

@[typedef]
pub struct C.VkVideoDecodeAV1CapabilitiesKHR {
pub mut:
	sType    StructureType = StructureType.video_decode_av1_capabilities_khr
	pNext    voidptr       = unsafe { nil }
	maxLevel StdVideoAV1Level
}

// VideoDecodeAV1SessionParametersCreateInfoKHR extends VkVideoSessionParametersCreateInfoKHR
pub type VideoDecodeAV1SessionParametersCreateInfoKHR = C.VkVideoDecodeAV1SessionParametersCreateInfoKHR

@[typedef]
pub struct C.VkVideoDecodeAV1SessionParametersCreateInfoKHR {
pub mut:
	sType              StructureType = StructureType.video_decode_av1_session_parameters_create_info_khr
	pNext              voidptr       = unsafe { nil }
	pStdSequenceHeader &StdVideoAV1SequenceHeader
}

// VideoDecodeAV1PictureInfoKHR extends VkVideoDecodeInfoKHR
pub type VideoDecodeAV1PictureInfoKHR = C.VkVideoDecodeAV1PictureInfoKHR

@[typedef]
pub struct C.VkVideoDecodeAV1PictureInfoKHR {
pub mut:
	sType                    StructureType = StructureType.video_decode_av1_picture_info_khr
	pNext                    voidptr       = unsafe { nil }
	pStdPictureInfo          &StdVideoDecodeAV1PictureInfo
	referenceNameSlotIndices [max_video_av1_references_per_frame_khr]i32
	frameHeaderOffset        u32
	tileCount                u32
	pTileOffsets             &u32
	pTileSizes               &u32
}

// VideoDecodeAV1DpbSlotInfoKHR extends VkVideoReferenceSlotInfoKHR
pub type VideoDecodeAV1DpbSlotInfoKHR = C.VkVideoDecodeAV1DpbSlotInfoKHR

@[typedef]
pub struct C.VkVideoDecodeAV1DpbSlotInfoKHR {
pub mut:
	sType             StructureType = StructureType.video_decode_av1_dpb_slot_info_khr
	pNext             voidptr       = unsafe { nil }
	pStdReferenceInfo &StdVideoDecodeAV1ReferenceInfo
}

pub const khr_video_encode_av1_spec_version = 1
pub const khr_video_encode_av1_extension_name = c'VK_KHR_video_encode_av1'

pub enum VideoEncodeAV1PredictionModeKHR as u32 {
	intra_only              = 0
	single_reference        = 1
	unidirectional_compound = 2
	bidirectional_compound  = 3
	max_enum_khr            = max_int
}

pub enum VideoEncodeAV1RateControlGroupKHR as u32 {
	intra        = 0
	predictive   = 1
	bipredictive = 2
	max_enum_khr = max_int
}

pub enum VideoEncodeAV1CapabilityFlagBitsKHR as u32 {
	per_rate_control_group_min_max_q_index = u32(0x00000001)
	generate_obu_extension_header          = u32(0x00000002)
	primary_reference_cdf_only             = u32(0x00000004)
	frame_size_override                    = u32(0x00000008)
	motion_vector_scaling                  = u32(0x00000010)
	compound_prediction_intra_refresh      = u32(0x00000020)
	max_enum_khr                           = max_int
}
pub type VideoEncodeAV1CapabilityFlagsKHR = u32

pub enum VideoEncodeAV1StdFlagBitsKHR as u32 {
	uniform_tile_spacing_flag_set = u32(0x00000001)
	skip_mode_present_unset       = u32(0x00000002)
	primary_ref_frame             = u32(0x00000004)
	delta_q                       = u32(0x00000008)
	max_enum_khr                  = max_int
}
pub type VideoEncodeAV1StdFlagsKHR = u32

pub enum VideoEncodeAV1SuperblockSizeFlagBitsKHR as u32 {
	_64          = u32(0x00000001)
	_128         = u32(0x00000002)
	max_enum_khr = max_int
}
pub type VideoEncodeAV1SuperblockSizeFlagsKHR = u32

pub enum VideoEncodeAV1RateControlFlagBitsKHR as u32 {
	regular_gop                   = u32(0x00000001)
	temporal_layer_pattern_dyadic = u32(0x00000002)
	reference_pattern_flat        = u32(0x00000004)
	reference_pattern_dyadic      = u32(0x00000008)
	max_enum_khr                  = max_int
}
pub type VideoEncodeAV1RateControlFlagsKHR = u32

// PhysicalDeviceVideoEncodeAV1FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVideoEncodeAV1FeaturesKHR = C.VkPhysicalDeviceVideoEncodeAV1FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceVideoEncodeAV1FeaturesKHR {
pub mut:
	sType          StructureType = StructureType.physical_device_video_encode_av1_features_khr
	pNext          voidptr       = unsafe { nil }
	videoEncodeAV1 Bool32
}

// VideoEncodeAV1CapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoEncodeAV1CapabilitiesKHR = C.VkVideoEncodeAV1CapabilitiesKHR

@[typedef]
pub struct C.VkVideoEncodeAV1CapabilitiesKHR {
pub mut:
	sType                                         StructureType = StructureType.video_encode_av1_capabilities_khr
	pNext                                         voidptr       = unsafe { nil }
	flags                                         VideoEncodeAV1CapabilityFlagsKHR
	maxLevel                                      StdVideoAV1Level
	codedPictureAlignment                         Extent2D
	maxTiles                                      Extent2D
	minTileSize                                   Extent2D
	maxTileSize                                   Extent2D
	superblockSizes                               VideoEncodeAV1SuperblockSizeFlagsKHR
	maxSingleReferenceCount                       u32
	singleReferenceNameMask                       u32
	maxUnidirectionalCompoundReferenceCount       u32
	maxUnidirectionalCompoundGroup1ReferenceCount u32
	unidirectionalCompoundReferenceNameMask       u32
	maxBidirectionalCompoundReferenceCount        u32
	maxBidirectionalCompoundGroup1ReferenceCount  u32
	maxBidirectionalCompoundGroup2ReferenceCount  u32
	bidirectionalCompoundReferenceNameMask        u32
	maxTemporalLayerCount                         u32
	maxSpatialLayerCount                          u32
	maxOperatingPoints                            u32
	minQIndex                                     u32
	maxQIndex                                     u32
	prefersGopRemainingFrames                     Bool32
	requiresGopRemainingFrames                    Bool32
	stdSyntaxFlags                                VideoEncodeAV1StdFlagsKHR
}

pub type VideoEncodeAV1QIndexKHR = C.VkVideoEncodeAV1QIndexKHR

@[typedef]
pub struct C.VkVideoEncodeAV1QIndexKHR {
pub mut:
	intraQIndex        u32
	predictiveQIndex   u32
	bipredictiveQIndex u32
}

// VideoEncodeAV1QualityLevelPropertiesKHR extends VkVideoEncodeQualityLevelPropertiesKHR
pub type VideoEncodeAV1QualityLevelPropertiesKHR = C.VkVideoEncodeAV1QualityLevelPropertiesKHR

@[typedef]
pub struct C.VkVideoEncodeAV1QualityLevelPropertiesKHR {
pub mut:
	sType                                                  StructureType = StructureType.video_encode_av1_quality_level_properties_khr
	pNext                                                  voidptr       = unsafe { nil }
	preferredRateControlFlags                              VideoEncodeAV1RateControlFlagsKHR
	preferredGopFrameCount                                 u32
	preferredKeyFramePeriod                                u32
	preferredConsecutiveBipredictiveFrameCount             u32
	preferredTemporalLayerCount                            u32
	preferredConstantQIndex                                VideoEncodeAV1QIndexKHR
	preferredMaxSingleReferenceCount                       u32
	preferredSingleReferenceNameMask                       u32
	preferredMaxUnidirectionalCompoundReferenceCount       u32
	preferredMaxUnidirectionalCompoundGroup1ReferenceCount u32
	preferredUnidirectionalCompoundReferenceNameMask       u32
	preferredMaxBidirectionalCompoundReferenceCount        u32
	preferredMaxBidirectionalCompoundGroup1ReferenceCount  u32
	preferredMaxBidirectionalCompoundGroup2ReferenceCount  u32
	preferredBidirectionalCompoundReferenceNameMask        u32
}

// VideoEncodeAV1SessionCreateInfoKHR extends VkVideoSessionCreateInfoKHR
pub type VideoEncodeAV1SessionCreateInfoKHR = C.VkVideoEncodeAV1SessionCreateInfoKHR

@[typedef]
pub struct C.VkVideoEncodeAV1SessionCreateInfoKHR {
pub mut:
	sType       StructureType = StructureType.video_encode_av1_session_create_info_khr
	pNext       voidptr       = unsafe { nil }
	useMaxLevel Bool32
	maxLevel    StdVideoAV1Level
}

// VideoEncodeAV1SessionParametersCreateInfoKHR extends VkVideoSessionParametersCreateInfoKHR
pub type VideoEncodeAV1SessionParametersCreateInfoKHR = C.VkVideoEncodeAV1SessionParametersCreateInfoKHR

@[typedef]
pub struct C.VkVideoEncodeAV1SessionParametersCreateInfoKHR {
pub mut:
	sType                  StructureType = StructureType.video_encode_av1_session_parameters_create_info_khr
	pNext                  voidptr       = unsafe { nil }
	pStdSequenceHeader     &StdVideoAV1SequenceHeader
	pStdDecoderModelInfo   &StdVideoEncodeAV1DecoderModelInfo
	stdOperatingPointCount u32
	pStdOperatingPoints    &StdVideoEncodeAV1OperatingPointInfo
}

// VideoEncodeAV1PictureInfoKHR extends VkVideoEncodeInfoKHR
pub type VideoEncodeAV1PictureInfoKHR = C.VkVideoEncodeAV1PictureInfoKHR

@[typedef]
pub struct C.VkVideoEncodeAV1PictureInfoKHR {
pub mut:
	sType                      StructureType = StructureType.video_encode_av1_picture_info_khr
	pNext                      voidptr       = unsafe { nil }
	predictionMode             VideoEncodeAV1PredictionModeKHR
	rateControlGroup           VideoEncodeAV1RateControlGroupKHR
	constantQIndex             u32
	pStdPictureInfo            &StdVideoEncodeAV1PictureInfo
	referenceNameSlotIndices   [max_video_av1_references_per_frame_khr]i32
	primaryReferenceCdfOnly    Bool32
	generateObuExtensionHeader Bool32
}

// VideoEncodeAV1DpbSlotInfoKHR extends VkVideoReferenceSlotInfoKHR
pub type VideoEncodeAV1DpbSlotInfoKHR = C.VkVideoEncodeAV1DpbSlotInfoKHR

@[typedef]
pub struct C.VkVideoEncodeAV1DpbSlotInfoKHR {
pub mut:
	sType             StructureType = StructureType.video_encode_av1_dpb_slot_info_khr
	pNext             voidptr       = unsafe { nil }
	pStdReferenceInfo &StdVideoEncodeAV1ReferenceInfo
}

// VideoEncodeAV1ProfileInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub type VideoEncodeAV1ProfileInfoKHR = C.VkVideoEncodeAV1ProfileInfoKHR

@[typedef]
pub struct C.VkVideoEncodeAV1ProfileInfoKHR {
pub mut:
	sType      StructureType = StructureType.video_encode_av1_profile_info_khr
	pNext      voidptr       = unsafe { nil }
	stdProfile StdVideoAV1Profile
}

pub type VideoEncodeAV1FrameSizeKHR = C.VkVideoEncodeAV1FrameSizeKHR

@[typedef]
pub struct C.VkVideoEncodeAV1FrameSizeKHR {
pub mut:
	intraFrameSize        u32
	predictiveFrameSize   u32
	bipredictiveFrameSize u32
}

// VideoEncodeAV1GopRemainingFrameInfoKHR extends VkVideoBeginCodingInfoKHR
pub type VideoEncodeAV1GopRemainingFrameInfoKHR = C.VkVideoEncodeAV1GopRemainingFrameInfoKHR

@[typedef]
pub struct C.VkVideoEncodeAV1GopRemainingFrameInfoKHR {
pub mut:
	sType                    StructureType = StructureType.video_encode_av1_gop_remaining_frame_info_khr
	pNext                    voidptr       = unsafe { nil }
	useGopRemainingFrames    Bool32
	gopRemainingIntra        u32
	gopRemainingPredictive   u32
	gopRemainingBipredictive u32
}

// VideoEncodeAV1RateControlInfoKHR extends VkVideoCodingControlInfoKHR,VkVideoBeginCodingInfoKHR
pub type VideoEncodeAV1RateControlInfoKHR = C.VkVideoEncodeAV1RateControlInfoKHR

@[typedef]
pub struct C.VkVideoEncodeAV1RateControlInfoKHR {
pub mut:
	sType                             StructureType = StructureType.video_encode_av1_rate_control_info_khr
	pNext                             voidptr       = unsafe { nil }
	flags                             VideoEncodeAV1RateControlFlagsKHR
	gopFrameCount                     u32
	keyFramePeriod                    u32
	consecutiveBipredictiveFrameCount u32
	temporalLayerCount                u32
}

// VideoEncodeAV1RateControlLayerInfoKHR extends VkVideoEncodeRateControlLayerInfoKHR
pub type VideoEncodeAV1RateControlLayerInfoKHR = C.VkVideoEncodeAV1RateControlLayerInfoKHR

@[typedef]
pub struct C.VkVideoEncodeAV1RateControlLayerInfoKHR {
pub mut:
	sType           StructureType = StructureType.video_encode_av1_rate_control_layer_info_khr
	pNext           voidptr       = unsafe { nil }
	useMinQIndex    Bool32
	minQIndex       VideoEncodeAV1QIndexKHR
	useMaxQIndex    Bool32
	maxQIndex       VideoEncodeAV1QIndexKHR
	useMaxFrameSize Bool32
	maxFrameSize    VideoEncodeAV1FrameSizeKHR
}

pub const max_video_vp9_references_per_frame_khr = u32(3)
pub const khr_video_decode_vp9_spec_version = 1
pub const khr_video_decode_vp9_extension_name = c'VK_KHR_video_decode_vp9'
// PhysicalDeviceVideoDecodeVP9FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVideoDecodeVP9FeaturesKHR = C.VkPhysicalDeviceVideoDecodeVP9FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceVideoDecodeVP9FeaturesKHR {
pub mut:
	sType          StructureType = StructureType.physical_device_video_decode_vp9_features_khr
	pNext          voidptr       = unsafe { nil }
	videoDecodeVP9 Bool32
}

// VideoDecodeVP9ProfileInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub type VideoDecodeVP9ProfileInfoKHR = C.VkVideoDecodeVP9ProfileInfoKHR

@[typedef]
pub struct C.VkVideoDecodeVP9ProfileInfoKHR {
pub mut:
	sType      StructureType = StructureType.video_decode_vp9_profile_info_khr
	pNext      voidptr       = unsafe { nil }
	stdProfile StdVideoVP9Profile
}

// VideoDecodeVP9CapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoDecodeVP9CapabilitiesKHR = C.VkVideoDecodeVP9CapabilitiesKHR

@[typedef]
pub struct C.VkVideoDecodeVP9CapabilitiesKHR {
pub mut:
	sType    StructureType = StructureType.video_decode_vp9_capabilities_khr
	pNext    voidptr       = unsafe { nil }
	maxLevel StdVideoVP9Level
}

// VideoDecodeVP9PictureInfoKHR extends VkVideoDecodeInfoKHR
pub type VideoDecodeVP9PictureInfoKHR = C.VkVideoDecodeVP9PictureInfoKHR

@[typedef]
pub struct C.VkVideoDecodeVP9PictureInfoKHR {
pub mut:
	sType                    StructureType = StructureType.video_decode_vp9_picture_info_khr
	pNext                    voidptr       = unsafe { nil }
	pStdPictureInfo          &StdVideoDecodeVP9PictureInfo
	referenceNameSlotIndices [max_video_vp9_references_per_frame_khr]i32
	uncompressedHeaderOffset u32
	compressedHeaderOffset   u32
	tilesOffset              u32
}

pub const khr_video_maintenance_1_spec_version = 1
pub const khr_video_maintenance_1_extension_name = c'VK_KHR_video_maintenance1'
// PhysicalDeviceVideoMaintenance1FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVideoMaintenance1FeaturesKHR = C.VkPhysicalDeviceVideoMaintenance1FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceVideoMaintenance1FeaturesKHR {
pub mut:
	sType             StructureType = StructureType.physical_device_video_maintenance1_features_khr
	pNext             voidptr       = unsafe { nil }
	videoMaintenance1 Bool32
}

// VideoInlineQueryInfoKHR extends VkVideoDecodeInfoKHR,VkVideoEncodeInfoKHR
pub type VideoInlineQueryInfoKHR = C.VkVideoInlineQueryInfoKHR

@[typedef]
pub struct C.VkVideoInlineQueryInfoKHR {
pub mut:
	sType      StructureType = StructureType.video_inline_query_info_khr
	pNext      voidptr       = unsafe { nil }
	queryPool  QueryPool
	firstQuery u32
	queryCount u32
}

pub const khr_vertex_attribute_divisor_spec_version = 1
pub const khr_vertex_attribute_divisor_extension_name = c'VK_KHR_vertex_attribute_divisor'

pub type PhysicalDeviceVertexAttributeDivisorPropertiesKHR = C.VkPhysicalDeviceVertexAttributeDivisorProperties

pub type VertexInputBindingDivisorDescriptionKHR = C.VkVertexInputBindingDivisorDescription

pub type PipelineVertexInputDivisorStateCreateInfoKHR = C.VkPipelineVertexInputDivisorStateCreateInfo

pub type PhysicalDeviceVertexAttributeDivisorFeaturesKHR = C.VkPhysicalDeviceVertexAttributeDivisorFeatures

pub const khr_load_store_op_none_spec_version = 1
pub const khr_load_store_op_none_extension_name = c'VK_KHR_load_store_op_none'

pub const khr_unified_image_layouts_spec_version = 1
pub const khr_unified_image_layouts_extension_name = c'VK_KHR_unified_image_layouts'
// PhysicalDeviceUnifiedImageLayoutsFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceUnifiedImageLayoutsFeaturesKHR = C.VkPhysicalDeviceUnifiedImageLayoutsFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceUnifiedImageLayoutsFeaturesKHR {
pub mut:
	sType                    StructureType = StructureType.physical_device_unified_image_layouts_features_khr
	pNext                    voidptr       = unsafe { nil }
	unifiedImageLayouts      Bool32
	unifiedImageLayoutsVideo Bool32
}

// AttachmentFeedbackLoopInfoEXT extends VkRenderingAttachmentInfo
pub type AttachmentFeedbackLoopInfoEXT = C.VkAttachmentFeedbackLoopInfoEXT

@[typedef]
pub struct C.VkAttachmentFeedbackLoopInfoEXT {
pub mut:
	sType              StructureType = StructureType.attachment_feedback_loop_info_ext
	pNext              voidptr       = unsafe { nil }
	feedbackLoopEnable Bool32
}

pub const khr_shader_float_controls_2_spec_version = 1
pub const khr_shader_float_controls_2_extension_name = c'VK_KHR_shader_float_controls2'

pub type PhysicalDeviceShaderFloatControls2FeaturesKHR = C.VkPhysicalDeviceShaderFloatControls2Features

pub const khr_index_type_uint8_spec_version = 1
pub const khr_index_type_uint8_extension_name = c'VK_KHR_index_type_uint8'

pub type PhysicalDeviceIndexTypeUint8FeaturesKHR = C.VkPhysicalDeviceIndexTypeUint8Features

pub const khr_line_rasterization_spec_version = 1
pub const khr_line_rasterization_extension_name = c'VK_KHR_line_rasterization'

pub type LineRasterizationModeKHR = LineRasterizationMode

pub type PhysicalDeviceLineRasterizationFeaturesKHR = C.VkPhysicalDeviceLineRasterizationFeatures

pub type PhysicalDeviceLineRasterizationPropertiesKHR = C.VkPhysicalDeviceLineRasterizationProperties

pub type PipelineRasterizationLineStateCreateInfoKHR = C.VkPipelineRasterizationLineStateCreateInfo

@[keep_args_alive]
fn C.vkCmdSetLineStippleKHR(command_buffer CommandBuffer, line_stipple_factor u32, line_stipple_pattern u16)

pub type PFN_vkCmdSetLineStippleKHR = fn (command_buffer CommandBuffer, line_stipple_factor u32, line_stipple_pattern u16)

@[inline]
pub fn cmd_set_line_stipple_khr(command_buffer CommandBuffer,
	line_stipple_factor u32,
	line_stipple_pattern u16) {
	C.vkCmdSetLineStippleKHR(command_buffer, line_stipple_factor, line_stipple_pattern)
}

pub const khr_calibrated_timestamps_spec_version = 1
pub const khr_calibrated_timestamps_extension_name = c'VK_KHR_calibrated_timestamps'

pub enum TimeDomainKHR as u32 {
	device                    = 0
	clock_monotonic           = 1
	clock_monotonic_raw       = 2
	query_performance_counter = 3
	max_enum_khr              = max_int
}
pub type CalibratedTimestampInfoKHR = C.VkCalibratedTimestampInfoKHR

@[typedef]
pub struct C.VkCalibratedTimestampInfoKHR {
pub mut:
	sType      StructureType = StructureType.calibrated_timestamp_info_khr
	pNext      voidptr       = unsafe { nil }
	timeDomain TimeDomainKHR
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceCalibrateableTimeDomainsKHR(physical_device PhysicalDevice, p_time_domain_count &u32, p_time_domains &TimeDomainKHR) Result

pub type PFN_vkGetPhysicalDeviceCalibrateableTimeDomainsKHR = fn (physical_device PhysicalDevice, p_time_domain_count &u32, p_time_domains &TimeDomainKHR) Result

@[inline]
pub fn get_physical_device_calibrateable_time_domains_khr(physical_device PhysicalDevice,
	p_time_domain_count &u32,
	p_time_domains &TimeDomainKHR) Result {
	return C.vkGetPhysicalDeviceCalibrateableTimeDomainsKHR(physical_device, p_time_domain_count,
		p_time_domains)
}

@[keep_args_alive]
fn C.vkGetCalibratedTimestampsKHR(device Device, timestamp_count u32, p_timestamp_infos &CalibratedTimestampInfoKHR, p_timestamps &u64, p_max_deviation &u64) Result

pub type PFN_vkGetCalibratedTimestampsKHR = fn (device Device, timestamp_count u32, p_timestamp_infos &CalibratedTimestampInfoKHR, p_timestamps &u64, p_max_deviation &u64) Result

@[inline]
pub fn get_calibrated_timestamps_khr(device Device,
	timestamp_count u32,
	p_timestamp_infos &CalibratedTimestampInfoKHR,
	p_timestamps &u64,
	p_max_deviation &u64) Result {
	return C.vkGetCalibratedTimestampsKHR(device, timestamp_count, p_timestamp_infos,
		p_timestamps, p_max_deviation)
}

pub const khr_shader_expect_assume_spec_version = 1
pub const khr_shader_expect_assume_extension_name = c'VK_KHR_shader_expect_assume'

pub type PhysicalDeviceShaderExpectAssumeFeaturesKHR = C.VkPhysicalDeviceShaderExpectAssumeFeatures

pub const khr_maintenance_6_spec_version = 1
pub const khr_maintenance_6_extension_name = c'VK_KHR_maintenance6'

pub type PhysicalDeviceMaintenance6FeaturesKHR = C.VkPhysicalDeviceMaintenance6Features

pub type PhysicalDeviceMaintenance6PropertiesKHR = C.VkPhysicalDeviceMaintenance6Properties

pub type BindMemoryStatusKHR = C.VkBindMemoryStatus

pub type BindDescriptorSetsInfoKHR = C.VkBindDescriptorSetsInfo

pub type PushConstantsInfoKHR = C.VkPushConstantsInfo

pub type PushDescriptorSetInfoKHR = C.VkPushDescriptorSetInfo

pub type PushDescriptorSetWithTemplateInfoKHR = C.VkPushDescriptorSetWithTemplateInfo

pub type SetDescriptorBufferOffsetsInfoEXT = C.VkSetDescriptorBufferOffsetsInfoEXT

@[typedef]
pub struct C.VkSetDescriptorBufferOffsetsInfoEXT {
pub mut:
	sType          StructureType = StructureType.set_descriptor_buffer_offsets_info_ext
	pNext          voidptr       = unsafe { nil }
	stageFlags     ShaderStageFlags
	layout         PipelineLayout
	firstSet       u32
	setCount       u32
	pBufferIndices &u32
	pOffsets       &DeviceSize
}

pub type BindDescriptorBufferEmbeddedSamplersInfoEXT = C.VkBindDescriptorBufferEmbeddedSamplersInfoEXT

@[typedef]
pub struct C.VkBindDescriptorBufferEmbeddedSamplersInfoEXT {
pub mut:
	sType      StructureType = StructureType.bind_descriptor_buffer_embedded_samplers_info_ext
	pNext      voidptr       = unsafe { nil }
	stageFlags ShaderStageFlags
	layout     PipelineLayout
	set        u32
}

@[keep_args_alive]
fn C.vkCmdBindDescriptorSets2KHR(command_buffer CommandBuffer, p_bind_descriptor_sets_info &BindDescriptorSetsInfo)

pub type PFN_vkCmdBindDescriptorSets2KHR = fn (command_buffer CommandBuffer, p_bind_descriptor_sets_info &BindDescriptorSetsInfo)

@[inline]
pub fn cmd_bind_descriptor_sets2_khr(command_buffer CommandBuffer,
	p_bind_descriptor_sets_info &BindDescriptorSetsInfo) {
	C.vkCmdBindDescriptorSets2KHR(command_buffer, p_bind_descriptor_sets_info)
}

@[keep_args_alive]
fn C.vkCmdPushConstants2KHR(command_buffer CommandBuffer, p_push_constants_info &PushConstantsInfo)

pub type PFN_vkCmdPushConstants2KHR = fn (command_buffer CommandBuffer, p_push_constants_info &PushConstantsInfo)

@[inline]
pub fn cmd_push_constants2_khr(command_buffer CommandBuffer,
	p_push_constants_info &PushConstantsInfo) {
	C.vkCmdPushConstants2KHR(command_buffer, p_push_constants_info)
}

@[keep_args_alive]
fn C.vkCmdPushDescriptorSet2KHR(command_buffer CommandBuffer, p_push_descriptor_set_info &PushDescriptorSetInfo)

pub type PFN_vkCmdPushDescriptorSet2KHR = fn (command_buffer CommandBuffer, p_push_descriptor_set_info &PushDescriptorSetInfo)

@[inline]
pub fn cmd_push_descriptor_set2_khr(command_buffer CommandBuffer,
	p_push_descriptor_set_info &PushDescriptorSetInfo) {
	C.vkCmdPushDescriptorSet2KHR(command_buffer, p_push_descriptor_set_info)
}

@[keep_args_alive]
fn C.vkCmdPushDescriptorSetWithTemplate2KHR(command_buffer CommandBuffer, p_push_descriptor_set_with_template_info &PushDescriptorSetWithTemplateInfo)

pub type PFN_vkCmdPushDescriptorSetWithTemplate2KHR = fn (command_buffer CommandBuffer, p_push_descriptor_set_with_template_info &PushDescriptorSetWithTemplateInfo)

@[inline]
pub fn cmd_push_descriptor_set_with_template2_khr(command_buffer CommandBuffer,
	p_push_descriptor_set_with_template_info &PushDescriptorSetWithTemplateInfo) {
	C.vkCmdPushDescriptorSetWithTemplate2KHR(command_buffer, p_push_descriptor_set_with_template_info)
}

@[keep_args_alive]
fn C.vkCmdSetDescriptorBufferOffsets2EXT(command_buffer CommandBuffer, p_set_descriptor_buffer_offsets_info &SetDescriptorBufferOffsetsInfoEXT)

pub type PFN_vkCmdSetDescriptorBufferOffsets2EXT = fn (command_buffer CommandBuffer, p_set_descriptor_buffer_offsets_info &SetDescriptorBufferOffsetsInfoEXT)

@[inline]
pub fn cmd_set_descriptor_buffer_offsets2_ext(command_buffer CommandBuffer,
	p_set_descriptor_buffer_offsets_info &SetDescriptorBufferOffsetsInfoEXT) {
	C.vkCmdSetDescriptorBufferOffsets2EXT(command_buffer, p_set_descriptor_buffer_offsets_info)
}

@[keep_args_alive]
fn C.vkCmdBindDescriptorBufferEmbeddedSamplers2EXT(command_buffer CommandBuffer, p_bind_descriptor_buffer_embedded_samplers_info &BindDescriptorBufferEmbeddedSamplersInfoEXT)

pub type PFN_vkCmdBindDescriptorBufferEmbeddedSamplers2EXT = fn (command_buffer CommandBuffer, p_bind_descriptor_buffer_embedded_samplers_info &BindDescriptorBufferEmbeddedSamplersInfoEXT)

@[inline]
pub fn cmd_bind_descriptor_buffer_embedded_samplers2_ext(command_buffer CommandBuffer,
	p_bind_descriptor_buffer_embedded_samplers_info &BindDescriptorBufferEmbeddedSamplersInfoEXT) {
	C.vkCmdBindDescriptorBufferEmbeddedSamplers2EXT(command_buffer, p_bind_descriptor_buffer_embedded_samplers_info)
}

pub const khr_copy_memory_indirect_spec_version = 1
pub const khr_copy_memory_indirect_extension_name = c'VK_KHR_copy_memory_indirect'

pub enum AddressCopyFlagBitsKHR as u32 {
	device_local = u32(0x00000001)
	sparse       = u32(0x00000002)
	protected    = u32(0x00000004)
	max_enum_khr = max_int
}
pub type AddressCopyFlagsKHR = u32
pub type StridedDeviceAddressRangeKHR = C.VkStridedDeviceAddressRangeKHR

@[typedef]
pub struct C.VkStridedDeviceAddressRangeKHR {
pub mut:
	address DeviceAddress
	size    DeviceSize
	stride  DeviceSize
}

pub type CopyMemoryIndirectCommandKHR = C.VkCopyMemoryIndirectCommandKHR

@[typedef]
pub struct C.VkCopyMemoryIndirectCommandKHR {
pub mut:
	srcAddress DeviceAddress
	dstAddress DeviceAddress
	size       DeviceSize
}

pub type CopyMemoryIndirectInfoKHR = C.VkCopyMemoryIndirectInfoKHR

@[typedef]
pub struct C.VkCopyMemoryIndirectInfoKHR {
pub mut:
	sType            StructureType = StructureType.copy_memory_indirect_info_khr
	pNext            voidptr       = unsafe { nil }
	srcCopyFlags     AddressCopyFlagsKHR
	dstCopyFlags     AddressCopyFlagsKHR
	copyCount        u32
	copyAddressRange StridedDeviceAddressRangeKHR
}

pub type CopyMemoryToImageIndirectCommandKHR = C.VkCopyMemoryToImageIndirectCommandKHR

@[typedef]
pub struct C.VkCopyMemoryToImageIndirectCommandKHR {
pub mut:
	srcAddress        DeviceAddress
	bufferRowLength   u32
	bufferImageHeight u32
	imageSubresource  ImageSubresourceLayers
	imageOffset       Offset3D
	imageExtent       Extent3D
}

pub type CopyMemoryToImageIndirectInfoKHR = C.VkCopyMemoryToImageIndirectInfoKHR

@[typedef]
pub struct C.VkCopyMemoryToImageIndirectInfoKHR {
pub mut:
	sType              StructureType = StructureType.copy_memory_to_image_indirect_info_khr
	pNext              voidptr       = unsafe { nil }
	srcCopyFlags       AddressCopyFlagsKHR
	copyCount          u32
	copyAddressRange   StridedDeviceAddressRangeKHR
	dstImage           Image
	dstImageLayout     ImageLayout
	pImageSubresources &ImageSubresourceLayers
}

// PhysicalDeviceCopyMemoryIndirectFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCopyMemoryIndirectFeaturesKHR = C.VkPhysicalDeviceCopyMemoryIndirectFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceCopyMemoryIndirectFeaturesKHR {
pub mut:
	sType                     StructureType = StructureType.physical_device_copy_memory_indirect_features_khr
	pNext                     voidptr       = unsafe { nil }
	indirectMemoryCopy        Bool32
	indirectMemoryToImageCopy Bool32
}

// PhysicalDeviceCopyMemoryIndirectPropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceCopyMemoryIndirectPropertiesKHR = C.VkPhysicalDeviceCopyMemoryIndirectPropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceCopyMemoryIndirectPropertiesKHR {
pub mut:
	sType           StructureType = StructureType.physical_device_copy_memory_indirect_properties_khr
	pNext           voidptr       = unsafe { nil }
	supportedQueues QueueFlags
}

@[keep_args_alive]
fn C.vkCmdCopyMemoryIndirectKHR(command_buffer CommandBuffer, p_copy_memory_indirect_info &CopyMemoryIndirectInfoKHR)

pub type PFN_vkCmdCopyMemoryIndirectKHR = fn (command_buffer CommandBuffer, p_copy_memory_indirect_info &CopyMemoryIndirectInfoKHR)

@[inline]
pub fn cmd_copy_memory_indirect_khr(command_buffer CommandBuffer,
	p_copy_memory_indirect_info &CopyMemoryIndirectInfoKHR) {
	C.vkCmdCopyMemoryIndirectKHR(command_buffer, p_copy_memory_indirect_info)
}

@[keep_args_alive]
fn C.vkCmdCopyMemoryToImageIndirectKHR(command_buffer CommandBuffer, p_copy_memory_to_image_indirect_info &CopyMemoryToImageIndirectInfoKHR)

pub type PFN_vkCmdCopyMemoryToImageIndirectKHR = fn (command_buffer CommandBuffer, p_copy_memory_to_image_indirect_info &CopyMemoryToImageIndirectInfoKHR)

@[inline]
pub fn cmd_copy_memory_to_image_indirect_khr(command_buffer CommandBuffer,
	p_copy_memory_to_image_indirect_info &CopyMemoryToImageIndirectInfoKHR) {
	C.vkCmdCopyMemoryToImageIndirectKHR(command_buffer, p_copy_memory_to_image_indirect_info)
}

pub const khr_video_encode_intra_refresh_spec_version = 1
pub const khr_video_encode_intra_refresh_extension_name = c'VK_KHR_video_encode_intra_refresh'

pub enum VideoEncodeIntraRefreshModeFlagBitsKHR as u32 {
	none                  = 0
	per_picture_partition = u32(0x00000001)
	block_based           = u32(0x00000002)
	block_row_based       = u32(0x00000004)
	block_column_based    = u32(0x00000008)
	max_enum_khr          = max_int
}
pub type VideoEncodeIntraRefreshModeFlagsKHR = u32

// VideoEncodeIntraRefreshCapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoEncodeIntraRefreshCapabilitiesKHR = C.VkVideoEncodeIntraRefreshCapabilitiesKHR

@[typedef]
pub struct C.VkVideoEncodeIntraRefreshCapabilitiesKHR {
pub mut:
	sType                                   StructureType = StructureType.video_encode_intra_refresh_capabilities_khr
	pNext                                   voidptr       = unsafe { nil }
	intraRefreshModes                       VideoEncodeIntraRefreshModeFlagsKHR
	maxIntraRefreshCycleDuration            u32
	maxIntraRefreshActiveReferencePictures  u32
	partitionIndependentIntraRefreshRegions Bool32
	nonRectangularIntraRefreshRegions       Bool32
}

// VideoEncodeSessionIntraRefreshCreateInfoKHR extends VkVideoSessionCreateInfoKHR
pub type VideoEncodeSessionIntraRefreshCreateInfoKHR = C.VkVideoEncodeSessionIntraRefreshCreateInfoKHR

@[typedef]
pub struct C.VkVideoEncodeSessionIntraRefreshCreateInfoKHR {
pub mut:
	sType            StructureType = StructureType.video_encode_session_intra_refresh_create_info_khr
	pNext            voidptr       = unsafe { nil }
	intraRefreshMode VideoEncodeIntraRefreshModeFlagBitsKHR
}

// VideoEncodeIntraRefreshInfoKHR extends VkVideoEncodeInfoKHR
pub type VideoEncodeIntraRefreshInfoKHR = C.VkVideoEncodeIntraRefreshInfoKHR

@[typedef]
pub struct C.VkVideoEncodeIntraRefreshInfoKHR {
pub mut:
	sType                     StructureType = StructureType.video_encode_intra_refresh_info_khr
	pNext                     voidptr       = unsafe { nil }
	intraRefreshCycleDuration u32
	intraRefreshIndex         u32
}

// VideoReferenceIntraRefreshInfoKHR extends VkVideoReferenceSlotInfoKHR
pub type VideoReferenceIntraRefreshInfoKHR = C.VkVideoReferenceIntraRefreshInfoKHR

@[typedef]
pub struct C.VkVideoReferenceIntraRefreshInfoKHR {
pub mut:
	sType                    StructureType = StructureType.video_reference_intra_refresh_info_khr
	pNext                    voidptr       = unsafe { nil }
	dirtyIntraRefreshRegions u32
}

// PhysicalDeviceVideoEncodeIntraRefreshFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVideoEncodeIntraRefreshFeaturesKHR = C.VkPhysicalDeviceVideoEncodeIntraRefreshFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceVideoEncodeIntraRefreshFeaturesKHR {
pub mut:
	sType                   StructureType = StructureType.physical_device_video_encode_intra_refresh_features_khr
	pNext                   voidptr       = unsafe { nil }
	videoEncodeIntraRefresh Bool32
}

pub const khr_video_encode_quantization_map_spec_version = 2
pub const khr_video_encode_quantization_map_extension_name = c'VK_KHR_video_encode_quantization_map'
// VideoEncodeQuantizationMapCapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoEncodeQuantizationMapCapabilitiesKHR = C.VkVideoEncodeQuantizationMapCapabilitiesKHR

@[typedef]
pub struct C.VkVideoEncodeQuantizationMapCapabilitiesKHR {
pub mut:
	sType                    StructureType = StructureType.video_encode_quantization_map_capabilities_khr
	pNext                    voidptr       = unsafe { nil }
	maxQuantizationMapExtent Extent2D
}

// VideoFormatQuantizationMapPropertiesKHR extends VkVideoFormatPropertiesKHR
pub type VideoFormatQuantizationMapPropertiesKHR = C.VkVideoFormatQuantizationMapPropertiesKHR

@[typedef]
pub struct C.VkVideoFormatQuantizationMapPropertiesKHR {
pub mut:
	sType                    StructureType = StructureType.video_format_quantization_map_properties_khr
	pNext                    voidptr       = unsafe { nil }
	quantizationMapTexelSize Extent2D
}

// VideoEncodeQuantizationMapInfoKHR extends VkVideoEncodeInfoKHR
pub type VideoEncodeQuantizationMapInfoKHR = C.VkVideoEncodeQuantizationMapInfoKHR

@[typedef]
pub struct C.VkVideoEncodeQuantizationMapInfoKHR {
pub mut:
	sType                 StructureType = StructureType.video_encode_quantization_map_info_khr
	pNext                 voidptr       = unsafe { nil }
	quantizationMap       ImageView
	quantizationMapExtent Extent2D
}

// VideoEncodeQuantizationMapSessionParametersCreateInfoKHR extends VkVideoSessionParametersCreateInfoKHR
pub type VideoEncodeQuantizationMapSessionParametersCreateInfoKHR = C.VkVideoEncodeQuantizationMapSessionParametersCreateInfoKHR

@[typedef]
pub struct C.VkVideoEncodeQuantizationMapSessionParametersCreateInfoKHR {
pub mut:
	sType                    StructureType = StructureType.video_encode_quantization_map_session_parameters_create_info_khr
	pNext                    voidptr       = unsafe { nil }
	quantizationMapTexelSize Extent2D
}

// PhysicalDeviceVideoEncodeQuantizationMapFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVideoEncodeQuantizationMapFeaturesKHR = C.VkPhysicalDeviceVideoEncodeQuantizationMapFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceVideoEncodeQuantizationMapFeaturesKHR {
pub mut:
	sType                      StructureType = StructureType.physical_device_video_encode_quantization_map_features_khr
	pNext                      voidptr       = unsafe { nil }
	videoEncodeQuantizationMap Bool32
}

// VideoEncodeH264QuantizationMapCapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoEncodeH264QuantizationMapCapabilitiesKHR = C.VkVideoEncodeH264QuantizationMapCapabilitiesKHR

@[typedef]
pub struct C.VkVideoEncodeH264QuantizationMapCapabilitiesKHR {
pub mut:
	sType      StructureType = StructureType.video_encode_h264_quantization_map_capabilities_khr
	pNext      voidptr       = unsafe { nil }
	minQpDelta i32
	maxQpDelta i32
}

// VideoEncodeH265QuantizationMapCapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoEncodeH265QuantizationMapCapabilitiesKHR = C.VkVideoEncodeH265QuantizationMapCapabilitiesKHR

@[typedef]
pub struct C.VkVideoEncodeH265QuantizationMapCapabilitiesKHR {
pub mut:
	sType      StructureType = StructureType.video_encode_h265_quantization_map_capabilities_khr
	pNext      voidptr       = unsafe { nil }
	minQpDelta i32
	maxQpDelta i32
}

// VideoFormatH265QuantizationMapPropertiesKHR extends VkVideoFormatPropertiesKHR
pub type VideoFormatH265QuantizationMapPropertiesKHR = C.VkVideoFormatH265QuantizationMapPropertiesKHR

@[typedef]
pub struct C.VkVideoFormatH265QuantizationMapPropertiesKHR {
pub mut:
	sType              StructureType = StructureType.video_format_h265_quantization_map_properties_khr
	pNext              voidptr       = unsafe { nil }
	compatibleCtbSizes VideoEncodeH265CtbSizeFlagsKHR
}

// VideoEncodeAV1QuantizationMapCapabilitiesKHR extends VkVideoCapabilitiesKHR
pub type VideoEncodeAV1QuantizationMapCapabilitiesKHR = C.VkVideoEncodeAV1QuantizationMapCapabilitiesKHR

@[typedef]
pub struct C.VkVideoEncodeAV1QuantizationMapCapabilitiesKHR {
pub mut:
	sType          StructureType = StructureType.video_encode_av1_quantization_map_capabilities_khr
	pNext          voidptr       = unsafe { nil }
	minQIndexDelta i32
	maxQIndexDelta i32
}

// VideoFormatAV1QuantizationMapPropertiesKHR extends VkVideoFormatPropertiesKHR
pub type VideoFormatAV1QuantizationMapPropertiesKHR = C.VkVideoFormatAV1QuantizationMapPropertiesKHR

@[typedef]
pub struct C.VkVideoFormatAV1QuantizationMapPropertiesKHR {
pub mut:
	sType                     StructureType = StructureType.video_format_av1_quantization_map_properties_khr
	pNext                     voidptr       = unsafe { nil }
	compatibleSuperblockSizes VideoEncodeAV1SuperblockSizeFlagsKHR
}

pub const khr_shader_relaxed_extended_instruction_spec_version = 1
pub const khr_shader_relaxed_extended_instruction_extension_name = c'VK_KHR_shader_relaxed_extended_instruction'
// PhysicalDeviceShaderRelaxedExtendedInstructionFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderRelaxedExtendedInstructionFeaturesKHR = C.VkPhysicalDeviceShaderRelaxedExtendedInstructionFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceShaderRelaxedExtendedInstructionFeaturesKHR {
pub mut:
	sType                            StructureType = StructureType.physical_device_shader_relaxed_extended_instruction_features_khr
	pNext                            voidptr       = unsafe { nil }
	shaderRelaxedExtendedInstruction Bool32
}

pub const khr_maintenance_7_spec_version = 1
pub const khr_maintenance_7_extension_name = c'VK_KHR_maintenance7'

pub enum PhysicalDeviceLayeredApiKHR as u32 {
	vulkan       = 0
	d3d12        = 1
	metal        = 2
	opengl       = 3
	opengles     = 4
	max_enum_khr = max_int
}
// PhysicalDeviceMaintenance7FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMaintenance7FeaturesKHR = C.VkPhysicalDeviceMaintenance7FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance7FeaturesKHR {
pub mut:
	sType        StructureType = StructureType.physical_device_maintenance7_features_khr
	pNext        voidptr       = unsafe { nil }
	maintenance7 Bool32
}

// PhysicalDeviceMaintenance7PropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMaintenance7PropertiesKHR = C.VkPhysicalDeviceMaintenance7PropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance7PropertiesKHR {
pub mut:
	sType                                                     StructureType = StructureType.physical_device_maintenance7_properties_khr
	pNext                                                     voidptr       = unsafe { nil }
	robustFragmentShadingRateAttachmentAccess                 Bool32
	separateDepthStencilAttachmentAccess                      Bool32
	maxDescriptorSetTotalUniformBuffersDynamic                u32
	maxDescriptorSetTotalStorageBuffersDynamic                u32
	maxDescriptorSetTotalBuffersDynamic                       u32
	maxDescriptorSetUpdateAfterBindTotalUniformBuffersDynamic u32
	maxDescriptorSetUpdateAfterBindTotalStorageBuffersDynamic u32
	maxDescriptorSetUpdateAfterBindTotalBuffersDynamic        u32
}

pub type PhysicalDeviceLayeredApiPropertiesKHR = C.VkPhysicalDeviceLayeredApiPropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceLayeredApiPropertiesKHR {
pub mut:
	sType      StructureType = StructureType.physical_device_layered_api_properties_khr
	pNext      voidptr       = unsafe { nil }
	vendorID   u32
	deviceID   u32
	layeredAPI PhysicalDeviceLayeredApiKHR
	deviceName [max_physical_device_name_size]char
}

// PhysicalDeviceLayeredApiPropertiesListKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceLayeredApiPropertiesListKHR = C.VkPhysicalDeviceLayeredApiPropertiesListKHR

@[typedef]
pub struct C.VkPhysicalDeviceLayeredApiPropertiesListKHR {
pub mut:
	sType           StructureType = StructureType.physical_device_layered_api_properties_list_khr
	pNext           voidptr       = unsafe { nil }
	layeredApiCount u32
	pLayeredApis    &PhysicalDeviceLayeredApiPropertiesKHR
}

// PhysicalDeviceLayeredApiVulkanPropertiesKHR extends VkPhysicalDeviceLayeredApiPropertiesKHR
pub type PhysicalDeviceLayeredApiVulkanPropertiesKHR = C.VkPhysicalDeviceLayeredApiVulkanPropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceLayeredApiVulkanPropertiesKHR {
pub mut:
	sType      StructureType = StructureType.physical_device_layered_api_vulkan_properties_khr
	pNext      voidptr       = unsafe { nil }
	properties PhysicalDeviceProperties2
}

pub const khr_maintenance_8_spec_version = 1
pub const khr_maintenance_8_extension_name = c'VK_KHR_maintenance8'

pub type AccessFlags3KHR = u64

// Flag bits for AccessFlagBits3KHR
pub type AccessFlagBits3KHR = u64

pub const access_3_none_khr = u64(0)

// MemoryBarrierAccessFlags3KHR extends VkSubpassDependency2,VkBufferMemoryBarrier2,VkImageMemoryBarrier2
pub type MemoryBarrierAccessFlags3KHR = C.VkMemoryBarrierAccessFlags3KHR

@[typedef]
pub struct C.VkMemoryBarrierAccessFlags3KHR {
pub mut:
	sType          StructureType = StructureType.memory_barrier_access_flags3_khr
	pNext          voidptr       = unsafe { nil }
	srcAccessMask3 AccessFlags3KHR
	dstAccessMask3 AccessFlags3KHR
}

// PhysicalDeviceMaintenance8FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMaintenance8FeaturesKHR = C.VkPhysicalDeviceMaintenance8FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance8FeaturesKHR {
pub mut:
	sType        StructureType = StructureType.physical_device_maintenance8_features_khr
	pNext        voidptr       = unsafe { nil }
	maintenance8 Bool32
}

pub const khr_shader_fma_spec_version = 1
pub const khr_shader_fma_extension_name = c'VK_KHR_shader_fma'
// PhysicalDeviceShaderFmaFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderFmaFeaturesKHR = C.VkPhysicalDeviceShaderFmaFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceShaderFmaFeaturesKHR {
pub mut:
	sType            StructureType = StructureType.physical_device_shader_fma_features_khr
	pNext            voidptr       = unsafe { nil }
	shaderFmaFloat16 Bool32
	shaderFmaFloat32 Bool32
	shaderFmaFloat64 Bool32
}

pub const khr_maintenance_9_spec_version = 1
pub const khr_maintenance_9_extension_name = c'VK_KHR_maintenance9'

pub enum DefaultVertexAttributeValueKHR as u32 {
	zero_zero_zero_zero = 0
	zero_zero_zero_one  = 1
	max_enum_khr        = max_int
}
// PhysicalDeviceMaintenance9FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMaintenance9FeaturesKHR = C.VkPhysicalDeviceMaintenance9FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance9FeaturesKHR {
pub mut:
	sType        StructureType = StructureType.physical_device_maintenance9_features_khr
	pNext        voidptr       = unsafe { nil }
	maintenance9 Bool32
}

// PhysicalDeviceMaintenance9PropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMaintenance9PropertiesKHR = C.VkPhysicalDeviceMaintenance9PropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance9PropertiesKHR {
pub mut:
	sType                       StructureType = StructureType.physical_device_maintenance9_properties_khr
	pNext                       voidptr       = unsafe { nil }
	image2DViewOf3DSparse       Bool32
	defaultVertexAttributeValue DefaultVertexAttributeValueKHR
}

// QueueFamilyOwnershipTransferPropertiesKHR extends VkQueueFamilyProperties2
pub type QueueFamilyOwnershipTransferPropertiesKHR = C.VkQueueFamilyOwnershipTransferPropertiesKHR

@[typedef]
pub struct C.VkQueueFamilyOwnershipTransferPropertiesKHR {
pub mut:
	sType                               StructureType = StructureType.queue_family_ownership_transfer_properties_khr
	pNext                               voidptr       = unsafe { nil }
	optimalImageTransferToQueueFamilies u32
}

pub const khr_video_maintenance_2_spec_version = 1
pub const khr_video_maintenance_2_extension_name = c'VK_KHR_video_maintenance2'
// PhysicalDeviceVideoMaintenance2FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVideoMaintenance2FeaturesKHR = C.VkPhysicalDeviceVideoMaintenance2FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceVideoMaintenance2FeaturesKHR {
pub mut:
	sType             StructureType = StructureType.physical_device_video_maintenance2_features_khr
	pNext             voidptr       = unsafe { nil }
	videoMaintenance2 Bool32
}

// VideoDecodeH264InlineSessionParametersInfoKHR extends VkVideoDecodeInfoKHR
pub type VideoDecodeH264InlineSessionParametersInfoKHR = C.VkVideoDecodeH264InlineSessionParametersInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH264InlineSessionParametersInfoKHR {
pub mut:
	sType   StructureType = StructureType.video_decode_h264_inline_session_parameters_info_khr
	pNext   voidptr       = unsafe { nil }
	pStdSPS &StdVideoH264SequenceParameterSet
	pStdPPS &StdVideoH264PictureParameterSet
}

// VideoDecodeH265InlineSessionParametersInfoKHR extends VkVideoDecodeInfoKHR
pub type VideoDecodeH265InlineSessionParametersInfoKHR = C.VkVideoDecodeH265InlineSessionParametersInfoKHR

@[typedef]
pub struct C.VkVideoDecodeH265InlineSessionParametersInfoKHR {
pub mut:
	sType   StructureType = StructureType.video_decode_h265_inline_session_parameters_info_khr
	pNext   voidptr       = unsafe { nil }
	pStdVPS &StdVideoH265VideoParameterSet
	pStdSPS &StdVideoH265SequenceParameterSet
	pStdPPS &StdVideoH265PictureParameterSet
}

// VideoDecodeAV1InlineSessionParametersInfoKHR extends VkVideoDecodeInfoKHR
pub type VideoDecodeAV1InlineSessionParametersInfoKHR = C.VkVideoDecodeAV1InlineSessionParametersInfoKHR

@[typedef]
pub struct C.VkVideoDecodeAV1InlineSessionParametersInfoKHR {
pub mut:
	sType              StructureType = StructureType.video_decode_av1_inline_session_parameters_info_khr
	pNext              voidptr       = unsafe { nil }
	pStdSequenceHeader &StdVideoAV1SequenceHeader
}

pub const khr_depth_clamp_zero_one_spec_version = 1
pub const khr_depth_clamp_zero_one_extension_name = c'VK_KHR_depth_clamp_zero_one'
// PhysicalDeviceDepthClampZeroOneFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDepthClampZeroOneFeaturesKHR = C.VkPhysicalDeviceDepthClampZeroOneFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceDepthClampZeroOneFeaturesKHR {
pub mut:
	sType             StructureType = StructureType.physical_device_depth_clamp_zero_one_features_khr
	pNext             voidptr       = unsafe { nil }
	depthClampZeroOne Bool32
}

pub const khr_robustness_2_spec_version = 1
pub const khr_robustness_2_extension_name = c'VK_KHR_robustness2'
// PhysicalDeviceRobustness2FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRobustness2FeaturesKHR = C.VkPhysicalDeviceRobustness2FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceRobustness2FeaturesKHR {
pub mut:
	sType               StructureType = StructureType.physical_device_robustness2_features_khr
	pNext               voidptr       = unsafe { nil }
	robustBufferAccess2 Bool32
	robustImageAccess2  Bool32
	nullDescriptor      Bool32
}

// PhysicalDeviceRobustness2PropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceRobustness2PropertiesKHR = C.VkPhysicalDeviceRobustness2PropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceRobustness2PropertiesKHR {
pub mut:
	sType                                  StructureType = StructureType.physical_device_robustness2_properties_khr
	pNext                                  voidptr       = unsafe { nil }
	robustStorageBufferAccessSizeAlignment DeviceSize
	robustUniformBufferAccessSizeAlignment DeviceSize
}

pub const khr_present_mode_fifo_latest_ready_spec_version = 1
pub const khr_present_mode_fifo_latest_ready_extension_name = c'VK_KHR_present_mode_fifo_latest_ready'
// PhysicalDevicePresentModeFifoLatestReadyFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePresentModeFifoLatestReadyFeaturesKHR = C.VkPhysicalDevicePresentModeFifoLatestReadyFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDevicePresentModeFifoLatestReadyFeaturesKHR {
pub mut:
	sType                      StructureType = StructureType.physical_device_present_mode_fifo_latest_ready_features_khr
	pNext                      voidptr       = unsafe { nil }
	presentModeFifoLatestReady Bool32
}

pub const khr_maintenance_10_spec_version = 1
pub const khr_maintenance_10_extension_name = c'VK_KHR_maintenance10'

pub enum RenderingAttachmentFlagBitsKHR as u32 {
	input_attachment_feedback        = u32(0x00000001)
	resolve_skip_transfer_function   = u32(0x00000002)
	resolve_enable_transfer_function = u32(0x00000004)
	max_enum_khr                     = max_int
}
pub type RenderingAttachmentFlagsKHR = u32

pub enum ResolveImageFlagBitsKHR as u32 {
	skip_transfer_function   = u32(0x00000001)
	enable_transfer_function = u32(0x00000002)
	max_enum_khr             = max_int
}
pub type ResolveImageFlagsKHR = u32

// PhysicalDeviceMaintenance10FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMaintenance10FeaturesKHR = C.VkPhysicalDeviceMaintenance10FeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance10FeaturesKHR {
pub mut:
	sType         StructureType = StructureType.physical_device_maintenance10_features_khr
	pNext         voidptr       = unsafe { nil }
	maintenance10 Bool32
}

// PhysicalDeviceMaintenance10PropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMaintenance10PropertiesKHR = C.VkPhysicalDeviceMaintenance10PropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceMaintenance10PropertiesKHR {
pub mut:
	sType                                            StructureType = StructureType.physical_device_maintenance10_properties_khr
	pNext                                            voidptr       = unsafe { nil }
	rgba4OpaqueBlackSwizzled                         Bool32
	resolveSrgbFormatAppliesTransferFunction         Bool32
	resolveSrgbFormatSupportsTransferFunctionControl Bool32
}

pub type RenderingEndInfoKHR = C.VkRenderingEndInfoKHR

@[typedef]
pub struct C.VkRenderingEndInfoKHR {
pub mut:
	sType StructureType = StructureType.rendering_end_info_khr
	pNext voidptr       = unsafe { nil }
}

// RenderingAttachmentFlagsInfoKHR extends VkRenderingAttachmentInfo
pub type RenderingAttachmentFlagsInfoKHR = C.VkRenderingAttachmentFlagsInfoKHR

@[typedef]
pub struct C.VkRenderingAttachmentFlagsInfoKHR {
pub mut:
	sType StructureType = StructureType.rendering_attachment_flags_info_khr
	pNext voidptr       = unsafe { nil }
	flags RenderingAttachmentFlagsKHR
}

// ResolveImageModeInfoKHR extends VkResolveImageInfo2
pub type ResolveImageModeInfoKHR = C.VkResolveImageModeInfoKHR

@[typedef]
pub struct C.VkResolveImageModeInfoKHR {
pub mut:
	sType              StructureType = StructureType.resolve_image_mode_info_khr
	pNext              voidptr       = unsafe { nil }
	flags              ResolveImageFlagsKHR
	resolveMode        ResolveModeFlagBits
	stencilResolveMode ResolveModeFlagBits
}

@[keep_args_alive]
fn C.vkCmdEndRendering2KHR(command_buffer CommandBuffer, p_rendering_end_info &RenderingEndInfoKHR)

pub type PFN_vkCmdEndRendering2KHR = fn (command_buffer CommandBuffer, p_rendering_end_info &RenderingEndInfoKHR)

@[inline]
pub fn cmd_end_rendering2_khr(command_buffer CommandBuffer,
	p_rendering_end_info &RenderingEndInfoKHR) {
	C.vkCmdEndRendering2KHR(command_buffer, p_rendering_end_info)
}

// Pointer to VkDebugReportCallbackEXT_T
pub type DebugReportCallbackEXT = voidptr

pub const ext_debug_report_spec_version = 10
pub const ext_debug_report_extension_name = c'VK_EXT_debug_report'

pub enum DebugReportObjectTypeEXT as u32 {
	unknown                    = 0
	instance                   = 1
	physical_device            = 2
	device                     = 3
	queue                      = 4
	semaphore                  = 5
	command_buffer             = 6
	fence                      = 7
	device_memory              = 8
	buffer                     = 9
	image                      = 10
	event                      = 11
	query_pool                 = 12
	buffer_view                = 13
	image_view                 = 14
	shader_module              = 15
	pipeline_cache             = 16
	pipeline_layout            = 17
	render_pass                = 18
	pipeline                   = 19
	descriptor_set_layout      = 20
	sampler                    = 21
	descriptor_pool            = 22
	descriptor_set             = 23
	framebuffer                = 24
	command_pool               = 25
	surface_khr                = 26
	swapchain_khr              = 27
	debug_report_callback_ext  = 28
	display_khr                = 29
	display_mode_khr           = 30
	validation_cache_ext       = 33
	sampler_ycbcr_conversion   = 1000156000
	descriptor_update_template = 1000085000
	cu_module_nvx              = 1000029000
	cu_function_nvx            = 1000029001
	acceleration_structure_khr = 1000150000
	acceleration_structure_nv  = 1000165000
	cuda_module_nv             = 1000307000
	cuda_function_nv           = 1000307001
	buffer_collection_fuchsia  = 1000366000
	max_enum_ext               = max_int
}

pub enum DebugReportFlagBitsEXT as u32 {
	information         = u32(0x00000001)
	warning             = u32(0x00000002)
	performance_warning = u32(0x00000004)
	error               = u32(0x00000008)
	debug               = u32(0x00000010)
	max_enum_ext        = max_int
}
pub type DebugReportFlagsEXT = u32
pub type PFN_vkDebugReportCallbackEXT = fn (DebugReportFlagsEXT, DebugReportObjectTypeEXT, u64, usize, i32, &char, &char, voidptr)

// DebugReportCallbackCreateInfoEXT extends VkInstanceCreateInfo
pub type DebugReportCallbackCreateInfoEXT = C.VkDebugReportCallbackCreateInfoEXT

@[typedef]
pub struct C.VkDebugReportCallbackCreateInfoEXT {
pub mut:
	sType       StructureType = StructureType.debug_report_callback_create_info_ext
	pNext       voidptr       = unsafe { nil }
	flags       DebugReportFlagsEXT
	pfnCallback PFN_vkDebugReportCallbackEXT = unsafe { nil }
	pUserData   voidptr                      = unsafe { nil }
}

@[keep_args_alive]
fn C.vkCreateDebugReportCallbackEXT(instance Instance, p_create_info &DebugReportCallbackCreateInfoEXT, p_allocator &AllocationCallbacks, p_callback &DebugReportCallbackEXT) Result

pub type PFN_vkCreateDebugReportCallbackEXT = fn (instance Instance, p_create_info &DebugReportCallbackCreateInfoEXT, p_allocator &AllocationCallbacks, p_callback &DebugReportCallbackEXT) Result

@[inline]
pub fn create_debug_report_callback_ext(instance Instance,
	p_create_info &DebugReportCallbackCreateInfoEXT,
	p_allocator &AllocationCallbacks,
	p_callback &DebugReportCallbackEXT) Result {
	return C.vkCreateDebugReportCallbackEXT(instance, p_create_info, p_allocator, p_callback)
}

@[keep_args_alive]
fn C.vkDestroyDebugReportCallbackEXT(instance Instance, callback DebugReportCallbackEXT, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyDebugReportCallbackEXT = fn (instance Instance, callback DebugReportCallbackEXT, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_debug_report_callback_ext(instance Instance,
	callback DebugReportCallbackEXT,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyDebugReportCallbackEXT(instance, callback, p_allocator)
}

@[keep_args_alive]
fn C.vkDebugReportMessageEXT(instance Instance, flags DebugReportFlagsEXT, object_type DebugReportObjectTypeEXT, object u64, location usize, message_code i32, p_layer_prefix &char, p_message &char)

pub type PFN_vkDebugReportMessageEXT = fn (instance Instance, flags DebugReportFlagsEXT, object_type DebugReportObjectTypeEXT, object u64, location usize, message_code i32, p_layer_prefix &char, p_message &char)

@[inline]
pub fn debug_report_message_ext(instance Instance,
	flags DebugReportFlagsEXT,
	object_type DebugReportObjectTypeEXT,
	object u64,
	location usize,
	message_code i32,
	p_layer_prefix &char,
	p_message &char) {
	C.vkDebugReportMessageEXT(instance, flags, object_type, object, location, message_code,
		p_layer_prefix, p_message)
}

pub const nv_glsl_shader_spec_version = 1
pub const nv_glsl_shader_extension_name = c'VK_NV_glsl_shader'

pub const ext_depth_range_unrestricted_spec_version = 1
pub const ext_depth_range_unrestricted_extension_name = c'VK_EXT_depth_range_unrestricted'

pub const img_filter_cubic_spec_version = 1
pub const img_filter_cubic_extension_name = c'VK_IMG_filter_cubic'

pub const amd_rasterization_order_spec_version = 1
pub const amd_rasterization_order_extension_name = c'VK_AMD_rasterization_order'

pub enum RasterizationOrderAMD as u32 {
	strict       = 0
	relaxed      = 1
	max_enum_amd = max_int
}
// PipelineRasterizationStateRasterizationOrderAMD extends VkPipelineRasterizationStateCreateInfo
pub type PipelineRasterizationStateRasterizationOrderAMD = C.VkPipelineRasterizationStateRasterizationOrderAMD

@[typedef]
pub struct C.VkPipelineRasterizationStateRasterizationOrderAMD {
pub mut:
	sType              StructureType = StructureType.pipeline_rasterization_state_rasterization_order_amd
	pNext              voidptr       = unsafe { nil }
	rasterizationOrder RasterizationOrderAMD
}

pub const amd_shader_trinary_minmax_spec_version = 1
pub const amd_shader_trinary_minmax_extension_name = c'VK_AMD_shader_trinary_minmax'

pub const amd_shader_explicit_vertex_parameter_spec_version = 1
pub const amd_shader_explicit_vertex_parameter_extension_name = c'VK_AMD_shader_explicit_vertex_parameter'

pub const ext_debug_marker_spec_version = 4
pub const ext_debug_marker_extension_name = c'VK_EXT_debug_marker'

pub type DebugMarkerObjectNameInfoEXT = C.VkDebugMarkerObjectNameInfoEXT

@[typedef]
pub struct C.VkDebugMarkerObjectNameInfoEXT {
pub mut:
	sType       StructureType = StructureType.debug_marker_object_name_info_ext
	pNext       voidptr       = unsafe { nil }
	objectType  DebugReportObjectTypeEXT
	object      u64
	pObjectName &char
}

pub type DebugMarkerObjectTagInfoEXT = C.VkDebugMarkerObjectTagInfoEXT

@[typedef]
pub struct C.VkDebugMarkerObjectTagInfoEXT {
pub mut:
	sType      StructureType = StructureType.debug_marker_object_tag_info_ext
	pNext      voidptr       = unsafe { nil }
	objectType DebugReportObjectTypeEXT
	object     u64
	tagName    u64
	tagSize    usize
	pTag       voidptr
}

pub type DebugMarkerMarkerInfoEXT = C.VkDebugMarkerMarkerInfoEXT

@[typedef]
pub struct C.VkDebugMarkerMarkerInfoEXT {
pub mut:
	sType       StructureType = StructureType.debug_marker_marker_info_ext
	pNext       voidptr       = unsafe { nil }
	pMarkerName &char
	color       [4]f32
}

@[keep_args_alive]
fn C.vkDebugMarkerSetObjectTagEXT(device Device, p_tag_info &DebugMarkerObjectTagInfoEXT) Result

pub type PFN_vkDebugMarkerSetObjectTagEXT = fn (device Device, p_tag_info &DebugMarkerObjectTagInfoEXT) Result

@[inline]
pub fn debug_marker_set_object_tag_ext(device Device,
	p_tag_info &DebugMarkerObjectTagInfoEXT) Result {
	return C.vkDebugMarkerSetObjectTagEXT(device, p_tag_info)
}

@[keep_args_alive]
fn C.vkDebugMarkerSetObjectNameEXT(device Device, p_name_info &DebugMarkerObjectNameInfoEXT) Result

pub type PFN_vkDebugMarkerSetObjectNameEXT = fn (device Device, p_name_info &DebugMarkerObjectNameInfoEXT) Result

@[inline]
pub fn debug_marker_set_object_name_ext(device Device,
	p_name_info &DebugMarkerObjectNameInfoEXT) Result {
	return C.vkDebugMarkerSetObjectNameEXT(device, p_name_info)
}

@[keep_args_alive]
fn C.vkCmdDebugMarkerBeginEXT(command_buffer CommandBuffer, p_marker_info &DebugMarkerMarkerInfoEXT)

pub type PFN_vkCmdDebugMarkerBeginEXT = fn (command_buffer CommandBuffer, p_marker_info &DebugMarkerMarkerInfoEXT)

@[inline]
pub fn cmd_debug_marker_begin_ext(command_buffer CommandBuffer,
	p_marker_info &DebugMarkerMarkerInfoEXT) {
	C.vkCmdDebugMarkerBeginEXT(command_buffer, p_marker_info)
}

@[keep_args_alive]
fn C.vkCmdDebugMarkerEndEXT(command_buffer CommandBuffer)

pub type PFN_vkCmdDebugMarkerEndEXT = fn (command_buffer CommandBuffer)

@[inline]
pub fn cmd_debug_marker_end_ext(command_buffer CommandBuffer) {
	C.vkCmdDebugMarkerEndEXT(command_buffer)
}

@[keep_args_alive]
fn C.vkCmdDebugMarkerInsertEXT(command_buffer CommandBuffer, p_marker_info &DebugMarkerMarkerInfoEXT)

pub type PFN_vkCmdDebugMarkerInsertEXT = fn (command_buffer CommandBuffer, p_marker_info &DebugMarkerMarkerInfoEXT)

@[inline]
pub fn cmd_debug_marker_insert_ext(command_buffer CommandBuffer,
	p_marker_info &DebugMarkerMarkerInfoEXT) {
	C.vkCmdDebugMarkerInsertEXT(command_buffer, p_marker_info)
}

pub const amd_gcn_shader_spec_version = 1
pub const amd_gcn_shader_extension_name = c'VK_AMD_gcn_shader'

pub const nv_dedicated_allocation_spec_version = 1
pub const nv_dedicated_allocation_extension_name = c'VK_NV_dedicated_allocation'
// DedicatedAllocationImageCreateInfoNV extends VkImageCreateInfo
pub type DedicatedAllocationImageCreateInfoNV = C.VkDedicatedAllocationImageCreateInfoNV

@[typedef]
pub struct C.VkDedicatedAllocationImageCreateInfoNV {
pub mut:
	sType               StructureType = StructureType.dedicated_allocation_image_create_info_nv
	pNext               voidptr       = unsafe { nil }
	dedicatedAllocation Bool32
}

// DedicatedAllocationBufferCreateInfoNV extends VkBufferCreateInfo
pub type DedicatedAllocationBufferCreateInfoNV = C.VkDedicatedAllocationBufferCreateInfoNV

@[typedef]
pub struct C.VkDedicatedAllocationBufferCreateInfoNV {
pub mut:
	sType               StructureType = StructureType.dedicated_allocation_buffer_create_info_nv
	pNext               voidptr       = unsafe { nil }
	dedicatedAllocation Bool32
}

// DedicatedAllocationMemoryAllocateInfoNV extends VkMemoryAllocateInfo
pub type DedicatedAllocationMemoryAllocateInfoNV = C.VkDedicatedAllocationMemoryAllocateInfoNV

@[typedef]
pub struct C.VkDedicatedAllocationMemoryAllocateInfoNV {
pub mut:
	sType  StructureType = StructureType.dedicated_allocation_memory_allocate_info_nv
	pNext  voidptr       = unsafe { nil }
	image  Image
	buffer Buffer
}

pub const ext_transform_feedback_spec_version = 1
pub const ext_transform_feedback_extension_name = c'VK_EXT_transform_feedback'

pub type PipelineRasterizationStateStreamCreateFlagsEXT = u32

// PhysicalDeviceTransformFeedbackFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceTransformFeedbackFeaturesEXT = C.VkPhysicalDeviceTransformFeedbackFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceTransformFeedbackFeaturesEXT {
pub mut:
	sType             StructureType = StructureType.physical_device_transform_feedback_features_ext
	pNext             voidptr       = unsafe { nil }
	transformFeedback Bool32
	geometryStreams   Bool32
}

// PhysicalDeviceTransformFeedbackPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceTransformFeedbackPropertiesEXT = C.VkPhysicalDeviceTransformFeedbackPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceTransformFeedbackPropertiesEXT {
pub mut:
	sType                                      StructureType = StructureType.physical_device_transform_feedback_properties_ext
	pNext                                      voidptr       = unsafe { nil }
	maxTransformFeedbackStreams                u32
	maxTransformFeedbackBuffers                u32
	maxTransformFeedbackBufferSize             DeviceSize
	maxTransformFeedbackStreamDataSize         u32
	maxTransformFeedbackBufferDataSize         u32
	maxTransformFeedbackBufferDataStride       u32
	transformFeedbackQueries                   Bool32
	transformFeedbackStreamsLinesTriangles     Bool32
	transformFeedbackRasterizationStreamSelect Bool32
	transformFeedbackDraw                      Bool32
}

// PipelineRasterizationStateStreamCreateInfoEXT extends VkPipelineRasterizationStateCreateInfo
pub type PipelineRasterizationStateStreamCreateInfoEXT = C.VkPipelineRasterizationStateStreamCreateInfoEXT

@[typedef]
pub struct C.VkPipelineRasterizationStateStreamCreateInfoEXT {
pub mut:
	sType               StructureType = StructureType.pipeline_rasterization_state_stream_create_info_ext
	pNext               voidptr       = unsafe { nil }
	flags               PipelineRasterizationStateStreamCreateFlagsEXT
	rasterizationStream u32
}

@[keep_args_alive]
fn C.vkCmdBindTransformFeedbackBuffersEXT(command_buffer CommandBuffer, first_binding u32, binding_count u32, p_buffers &Buffer, p_offsets &DeviceSize, p_sizes &DeviceSize)

pub type PFN_vkCmdBindTransformFeedbackBuffersEXT = fn (command_buffer CommandBuffer, first_binding u32, binding_count u32, p_buffers &Buffer, p_offsets &DeviceSize, p_sizes &DeviceSize)

@[inline]
pub fn cmd_bind_transform_feedback_buffers_ext(command_buffer CommandBuffer,
	first_binding u32,
	binding_count u32,
	p_buffers &Buffer,
	p_offsets &DeviceSize,
	p_sizes &DeviceSize) {
	C.vkCmdBindTransformFeedbackBuffersEXT(command_buffer, first_binding, binding_count,
		p_buffers, p_offsets, p_sizes)
}

@[keep_args_alive]
fn C.vkCmdBeginTransformFeedbackEXT(command_buffer CommandBuffer, first_counter_buffer u32, counter_buffer_count u32, p_counter_buffers &Buffer, p_counter_buffer_offsets &DeviceSize)

pub type PFN_vkCmdBeginTransformFeedbackEXT = fn (command_buffer CommandBuffer, first_counter_buffer u32, counter_buffer_count u32, p_counter_buffers &Buffer, p_counter_buffer_offsets &DeviceSize)

@[inline]
pub fn cmd_begin_transform_feedback_ext(command_buffer CommandBuffer,
	first_counter_buffer u32,
	counter_buffer_count u32,
	p_counter_buffers &Buffer,
	p_counter_buffer_offsets &DeviceSize) {
	C.vkCmdBeginTransformFeedbackEXT(command_buffer, first_counter_buffer, counter_buffer_count,
		p_counter_buffers, p_counter_buffer_offsets)
}

@[keep_args_alive]
fn C.vkCmdEndTransformFeedbackEXT(command_buffer CommandBuffer, first_counter_buffer u32, counter_buffer_count u32, p_counter_buffers &Buffer, p_counter_buffer_offsets &DeviceSize)

pub type PFN_vkCmdEndTransformFeedbackEXT = fn (command_buffer CommandBuffer, first_counter_buffer u32, counter_buffer_count u32, p_counter_buffers &Buffer, p_counter_buffer_offsets &DeviceSize)

@[inline]
pub fn cmd_end_transform_feedback_ext(command_buffer CommandBuffer,
	first_counter_buffer u32,
	counter_buffer_count u32,
	p_counter_buffers &Buffer,
	p_counter_buffer_offsets &DeviceSize) {
	C.vkCmdEndTransformFeedbackEXT(command_buffer, first_counter_buffer, counter_buffer_count,
		p_counter_buffers, p_counter_buffer_offsets)
}

@[keep_args_alive]
fn C.vkCmdBeginQueryIndexedEXT(command_buffer CommandBuffer, query_pool QueryPool, query u32, flags QueryControlFlags, index u32)

pub type PFN_vkCmdBeginQueryIndexedEXT = fn (command_buffer CommandBuffer, query_pool QueryPool, query u32, flags QueryControlFlags, index u32)

@[inline]
pub fn cmd_begin_query_indexed_ext(command_buffer CommandBuffer,
	query_pool QueryPool,
	query u32,
	flags QueryControlFlags,
	index u32) {
	C.vkCmdBeginQueryIndexedEXT(command_buffer, query_pool, query, flags, index)
}

@[keep_args_alive]
fn C.vkCmdEndQueryIndexedEXT(command_buffer CommandBuffer, query_pool QueryPool, query u32, index u32)

pub type PFN_vkCmdEndQueryIndexedEXT = fn (command_buffer CommandBuffer, query_pool QueryPool, query u32, index u32)

@[inline]
pub fn cmd_end_query_indexed_ext(command_buffer CommandBuffer,
	query_pool QueryPool,
	query u32,
	index u32) {
	C.vkCmdEndQueryIndexedEXT(command_buffer, query_pool, query, index)
}

@[keep_args_alive]
fn C.vkCmdDrawIndirectByteCountEXT(command_buffer CommandBuffer, instance_count u32, first_instance u32, counter_buffer Buffer, counter_buffer_offset DeviceSize, counter_offset u32, vertex_stride u32)

pub type PFN_vkCmdDrawIndirectByteCountEXT = fn (command_buffer CommandBuffer, instance_count u32, first_instance u32, counter_buffer Buffer, counter_buffer_offset DeviceSize, counter_offset u32, vertex_stride u32)

@[inline]
pub fn cmd_draw_indirect_byte_count_ext(command_buffer CommandBuffer,
	instance_count u32,
	first_instance u32,
	counter_buffer Buffer,
	counter_buffer_offset DeviceSize,
	counter_offset u32,
	vertex_stride u32) {
	C.vkCmdDrawIndirectByteCountEXT(command_buffer, instance_count, first_instance, counter_buffer,
		counter_buffer_offset, counter_offset, vertex_stride)
}

// Pointer to VkCuModuleNVX_T
pub type CuModuleNVX = voidptr

// Pointer to VkCuFunctionNVX_T
pub type CuFunctionNVX = voidptr

pub const nvx_binary_import_spec_version = 2
pub const nvx_binary_import_extension_name = c'VK_NVX_binary_import'

pub type CuModuleCreateInfoNVX = C.VkCuModuleCreateInfoNVX

@[typedef]
pub struct C.VkCuModuleCreateInfoNVX {
pub mut:
	sType    StructureType = StructureType.cu_module_create_info_nvx
	pNext    voidptr       = unsafe { nil }
	dataSize usize
	pData    voidptr
}

// CuModuleTexturingModeCreateInfoNVX extends VkCuModuleCreateInfoNVX
pub type CuModuleTexturingModeCreateInfoNVX = C.VkCuModuleTexturingModeCreateInfoNVX

@[typedef]
pub struct C.VkCuModuleTexturingModeCreateInfoNVX {
pub mut:
	sType             StructureType = StructureType.cu_module_texturing_mode_create_info_nvx
	pNext             voidptr       = unsafe { nil }
	use64bitTexturing Bool32
}

pub type CuFunctionCreateInfoNVX = C.VkCuFunctionCreateInfoNVX

@[typedef]
pub struct C.VkCuFunctionCreateInfoNVX {
pub mut:
	sType  StructureType = StructureType.cu_function_create_info_nvx
	pNext  voidptr       = unsafe { nil }
	module CuModuleNVX
	pName  &char
}

pub type CuLaunchInfoNVX = C.VkCuLaunchInfoNVX

@[typedef]
pub struct C.VkCuLaunchInfoNVX {
pub mut:
	sType          StructureType = StructureType.cu_launch_info_nvx
	pNext          voidptr       = unsafe { nil }
	function       CuFunctionNVX
	gridDimX       u32
	gridDimY       u32
	gridDimZ       u32
	blockDimX      u32
	blockDimY      u32
	blockDimZ      u32
	sharedMemBytes u32
	paramCount     usize
	pParams        &voidptr
	extraCount     usize
	pExtras        &voidptr
}

@[keep_args_alive]
fn C.vkCreateCuModuleNVX(device Device, p_create_info &CuModuleCreateInfoNVX, p_allocator &AllocationCallbacks, p_module &CuModuleNVX) Result

pub type PFN_vkCreateCuModuleNVX = fn (device Device, p_create_info &CuModuleCreateInfoNVX, p_allocator &AllocationCallbacks, p_module &CuModuleNVX) Result

@[inline]
pub fn create_cu_module_nvx(device Device,
	p_create_info &CuModuleCreateInfoNVX,
	p_allocator &AllocationCallbacks,
	p_module &CuModuleNVX) Result {
	return C.vkCreateCuModuleNVX(device, p_create_info, p_allocator, p_module)
}

@[keep_args_alive]
fn C.vkCreateCuFunctionNVX(device Device, p_create_info &CuFunctionCreateInfoNVX, p_allocator &AllocationCallbacks, p_function &CuFunctionNVX) Result

pub type PFN_vkCreateCuFunctionNVX = fn (device Device, p_create_info &CuFunctionCreateInfoNVX, p_allocator &AllocationCallbacks, p_function &CuFunctionNVX) Result

@[inline]
pub fn create_cu_function_nvx(device Device,
	p_create_info &CuFunctionCreateInfoNVX,
	p_allocator &AllocationCallbacks,
	p_function &CuFunctionNVX) Result {
	return C.vkCreateCuFunctionNVX(device, p_create_info, p_allocator, p_function)
}

@[keep_args_alive]
fn C.vkDestroyCuModuleNVX(device Device, vkmodule CuModuleNVX, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyCuModuleNVX = fn (device Device, vkmodule CuModuleNVX, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_cu_module_nvx(device Device,
	vkmodule CuModuleNVX,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyCuModuleNVX(device, vkmodule, p_allocator)
}

@[keep_args_alive]
fn C.vkDestroyCuFunctionNVX(device Device, function CuFunctionNVX, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyCuFunctionNVX = fn (device Device, function CuFunctionNVX, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_cu_function_nvx(device Device,
	function CuFunctionNVX,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyCuFunctionNVX(device, function, p_allocator)
}

@[keep_args_alive]
fn C.vkCmdCuLaunchKernelNVX(command_buffer CommandBuffer, p_launch_info &CuLaunchInfoNVX)

pub type PFN_vkCmdCuLaunchKernelNVX = fn (command_buffer CommandBuffer, p_launch_info &CuLaunchInfoNVX)

@[inline]
pub fn cmd_cu_launch_kernel_nvx(command_buffer CommandBuffer,
	p_launch_info &CuLaunchInfoNVX) {
	C.vkCmdCuLaunchKernelNVX(command_buffer, p_launch_info)
}

pub const nvx_image_view_handle_spec_version = 3
pub const nvx_image_view_handle_extension_name = c'VK_NVX_image_view_handle'

pub type ImageViewHandleInfoNVX = C.VkImageViewHandleInfoNVX

@[typedef]
pub struct C.VkImageViewHandleInfoNVX {
pub mut:
	sType          StructureType = StructureType.image_view_handle_info_nvx
	pNext          voidptr       = unsafe { nil }
	imageView      ImageView
	descriptorType DescriptorType
	sampler        Sampler
}

pub type ImageViewAddressPropertiesNVX = C.VkImageViewAddressPropertiesNVX

@[typedef]
pub struct C.VkImageViewAddressPropertiesNVX {
pub mut:
	sType         StructureType = StructureType.image_view_address_properties_nvx
	pNext         voidptr       = unsafe { nil }
	deviceAddress DeviceAddress
	size          DeviceSize
}

@[keep_args_alive]
fn C.vkGetImageViewHandleNVX(device Device, p_info &ImageViewHandleInfoNVX) u32

pub type PFN_vkGetImageViewHandleNVX = fn (device Device, p_info &ImageViewHandleInfoNVX) u32

@[inline]
pub fn get_image_view_handle_nvx(device Device,
	p_info &ImageViewHandleInfoNVX) u32 {
	return C.vkGetImageViewHandleNVX(device, p_info)
}

@[keep_args_alive]
fn C.vkGetImageViewHandle64NVX(device Device, p_info &ImageViewHandleInfoNVX) u64

pub type PFN_vkGetImageViewHandle64NVX = fn (device Device, p_info &ImageViewHandleInfoNVX) u64

@[inline]
pub fn get_image_view_handle64_nvx(device Device,
	p_info &ImageViewHandleInfoNVX) u64 {
	return C.vkGetImageViewHandle64NVX(device, p_info)
}

@[keep_args_alive]
fn C.vkGetImageViewAddressNVX(device Device, image_view ImageView, mut p_properties ImageViewAddressPropertiesNVX) Result

pub type PFN_vkGetImageViewAddressNVX = fn (device Device, image_view ImageView, mut p_properties ImageViewAddressPropertiesNVX) Result

@[inline]
pub fn get_image_view_address_nvx(device Device,
	image_view ImageView,
	mut p_properties ImageViewAddressPropertiesNVX) Result {
	return C.vkGetImageViewAddressNVX(device, image_view, mut p_properties)
}

pub const amd_draw_indirect_count_spec_version = 2
pub const amd_draw_indirect_count_extension_name = c'VK_AMD_draw_indirect_count'

@[keep_args_alive]
fn C.vkCmdDrawIndirectCountAMD(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

pub type PFN_vkCmdDrawIndirectCountAMD = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_indirect_count_amd(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	count_buffer Buffer,
	count_buffer_offset DeviceSize,
	max_draw_count u32,
	stride u32) {
	C.vkCmdDrawIndirectCountAMD(command_buffer, buffer, offset, count_buffer, count_buffer_offset,
		max_draw_count, stride)
}

@[keep_args_alive]
fn C.vkCmdDrawIndexedIndirectCountAMD(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

pub type PFN_vkCmdDrawIndexedIndirectCountAMD = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_indexed_indirect_count_amd(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	count_buffer Buffer,
	count_buffer_offset DeviceSize,
	max_draw_count u32,
	stride u32) {
	C.vkCmdDrawIndexedIndirectCountAMD(command_buffer, buffer, offset, count_buffer, count_buffer_offset,
		max_draw_count, stride)
}

pub const amd_negative_viewport_height_spec_version = 1
pub const amd_negative_viewport_height_extension_name = c'VK_AMD_negative_viewport_height'

pub const amd_gpu_shader_half_float_spec_version = 2
pub const amd_gpu_shader_half_float_extension_name = c'VK_AMD_gpu_shader_half_float'

pub const amd_shader_ballot_spec_version = 1
pub const amd_shader_ballot_extension_name = c'VK_AMD_shader_ballot'

pub const amd_texture_gather_bias_lod_spec_version = 1
pub const amd_texture_gather_bias_lod_extension_name = c'VK_AMD_texture_gather_bias_lod'
// TextureLODGatherFormatPropertiesAMD extends VkImageFormatProperties2
pub type TextureLODGatherFormatPropertiesAMD = C.VkTextureLODGatherFormatPropertiesAMD

@[typedef]
pub struct C.VkTextureLODGatherFormatPropertiesAMD {
pub mut:
	sType                           StructureType = StructureType.texture_lod_gather_format_properties_amd
	pNext                           voidptr       = unsafe { nil }
	supportsTextureGatherLODBiasAMD Bool32
}

pub const amd_shader_info_spec_version = 1
pub const amd_shader_info_extension_name = c'VK_AMD_shader_info'

pub enum ShaderInfoTypeAMD as u32 {
	statistics   = 0
	binary       = 1
	disassembly  = 2
	max_enum_amd = max_int
}
pub type ShaderResourceUsageAMD = C.VkShaderResourceUsageAMD

@[typedef]
pub struct C.VkShaderResourceUsageAMD {
pub mut:
	numUsedVgprs             u32
	numUsedSgprs             u32
	ldsSizePerLocalWorkGroup u32
	ldsUsageSizeInBytes      usize
	scratchMemUsageInBytes   usize
}

pub type ShaderStatisticsInfoAMD = C.VkShaderStatisticsInfoAMD

@[typedef]
pub struct C.VkShaderStatisticsInfoAMD {
pub mut:
	shaderStageMask      ShaderStageFlags
	resourceUsage        ShaderResourceUsageAMD
	numPhysicalVgprs     u32
	numPhysicalSgprs     u32
	numAvailableVgprs    u32
	numAvailableSgprs    u32
	computeWorkGroupSize [3]u32
}

@[keep_args_alive]
fn C.vkGetShaderInfoAMD(device Device, pipeline Pipeline, shader_stage ShaderStageFlagBits, info_type ShaderInfoTypeAMD, p_info_size &usize, p_info voidptr) Result

pub type PFN_vkGetShaderInfoAMD = fn (device Device, pipeline Pipeline, shader_stage ShaderStageFlagBits, info_type ShaderInfoTypeAMD, p_info_size &usize, p_info voidptr) Result

@[inline]
pub fn get_shader_info_amd(device Device,
	pipeline Pipeline,
	shader_stage ShaderStageFlagBits,
	info_type ShaderInfoTypeAMD,
	p_info_size &usize,
	p_info voidptr) Result {
	return C.vkGetShaderInfoAMD(device, pipeline, shader_stage, info_type, p_info_size,
		p_info)
}

pub const amd_shader_image_load_store_lod_spec_version = 1
pub const amd_shader_image_load_store_lod_extension_name = c'VK_AMD_shader_image_load_store_lod'

pub const nv_corner_sampled_image_spec_version = 2
pub const nv_corner_sampled_image_extension_name = c'VK_NV_corner_sampled_image'
// PhysicalDeviceCornerSampledImageFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCornerSampledImageFeaturesNV = C.VkPhysicalDeviceCornerSampledImageFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceCornerSampledImageFeaturesNV {
pub mut:
	sType              StructureType = StructureType.physical_device_corner_sampled_image_features_nv
	pNext              voidptr       = unsafe { nil }
	cornerSampledImage Bool32
}

pub const img_format_pvrtc_spec_version = 1
pub const img_format_pvrtc_extension_name = c'VK_IMG_format_pvrtc'

pub const nv_external_memory_capabilities_spec_version = 1
pub const nv_external_memory_capabilities_extension_name = c'VK_NV_external_memory_capabilities'

pub enum ExternalMemoryHandleTypeFlagBitsNV as u32 {
	opaque_win32     = u32(0x00000001)
	opaque_win32_kmt = u32(0x00000002)
	d3d11_image      = u32(0x00000004)
	d3d11_image_kmt  = u32(0x00000008)
	max_enum_nv      = max_int
}
pub type ExternalMemoryHandleTypeFlagsNV = u32

pub enum ExternalMemoryFeatureFlagBitsNV as u32 {
	dedicated_only = u32(0x00000001)
	exportable     = u32(0x00000002)
	importable     = u32(0x00000004)
	max_enum_nv    = max_int
}
pub type ExternalMemoryFeatureFlagsNV = u32
pub type ExternalImageFormatPropertiesNV = C.VkExternalImageFormatPropertiesNV

@[typedef]
pub struct C.VkExternalImageFormatPropertiesNV {
pub mut:
	imageFormatProperties         ImageFormatProperties
	externalMemoryFeatures        ExternalMemoryFeatureFlagsNV
	exportFromImportedHandleTypes ExternalMemoryHandleTypeFlagsNV
	compatibleHandleTypes         ExternalMemoryHandleTypeFlagsNV
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceExternalImageFormatPropertiesNV(physical_device PhysicalDevice, format Format, type_param ImageType, tiling ImageTiling, usage ImageUsageFlags, flags ImageCreateFlags, external_handle_type ExternalMemoryHandleTypeFlagsNV, mut p_external_image_format_properties ExternalImageFormatPropertiesNV) Result

pub type PFN_vkGetPhysicalDeviceExternalImageFormatPropertiesNV = fn (physical_device PhysicalDevice, format Format, type_param ImageType, tiling ImageTiling, usage ImageUsageFlags, flags ImageCreateFlags, external_handle_type ExternalMemoryHandleTypeFlagsNV, mut p_external_image_format_properties ExternalImageFormatPropertiesNV) Result

@[inline]
pub fn get_physical_device_external_image_format_properties_nv(physical_device PhysicalDevice,
	format Format,
	type_param ImageType,
	tiling ImageTiling,
	usage ImageUsageFlags,
	flags ImageCreateFlags,
	external_handle_type ExternalMemoryHandleTypeFlagsNV,
	mut p_external_image_format_properties ExternalImageFormatPropertiesNV) Result {
	return C.vkGetPhysicalDeviceExternalImageFormatPropertiesNV(physical_device, format,
		type_param, tiling, usage, flags, external_handle_type, mut p_external_image_format_properties)
}

pub const nv_external_memory_spec_version = 1
pub const nv_external_memory_extension_name = c'VK_NV_external_memory'
// ExternalMemoryImageCreateInfoNV extends VkImageCreateInfo
pub type ExternalMemoryImageCreateInfoNV = C.VkExternalMemoryImageCreateInfoNV

@[typedef]
pub struct C.VkExternalMemoryImageCreateInfoNV {
pub mut:
	sType       StructureType = StructureType.external_memory_image_create_info_nv
	pNext       voidptr       = unsafe { nil }
	handleTypes ExternalMemoryHandleTypeFlagsNV
}

// ExportMemoryAllocateInfoNV extends VkMemoryAllocateInfo
pub type ExportMemoryAllocateInfoNV = C.VkExportMemoryAllocateInfoNV

@[typedef]
pub struct C.VkExportMemoryAllocateInfoNV {
pub mut:
	sType       StructureType = StructureType.export_memory_allocate_info_nv
	pNext       voidptr       = unsafe { nil }
	handleTypes ExternalMemoryHandleTypeFlagsNV
}

pub const ext_validation_flags_spec_version = 3
pub const ext_validation_flags_extension_name = c'VK_EXT_validation_flags'

pub enum ValidationCheckEXT as u32 {
	all          = 0
	shaders      = 1
	max_enum_ext = max_int
}
// ValidationFlagsEXT extends VkInstanceCreateInfo
pub type ValidationFlagsEXT = C.VkValidationFlagsEXT

@[typedef]
pub struct C.VkValidationFlagsEXT {
pub mut:
	sType                        StructureType = StructureType.validation_flags_ext
	pNext                        voidptr       = unsafe { nil }
	disabledValidationCheckCount u32
	pDisabledValidationChecks    &ValidationCheckEXT
}

pub const ext_shader_subgroup_ballot_spec_version = 1
pub const ext_shader_subgroup_ballot_extension_name = c'VK_EXT_shader_subgroup_ballot'

pub const ext_shader_subgroup_vote_spec_version = 1
pub const ext_shader_subgroup_vote_extension_name = c'VK_EXT_shader_subgroup_vote'

pub const ext_texture_compression_astc_hdr_spec_version = 1
pub const ext_texture_compression_astc_hdr_extension_name = c'VK_EXT_texture_compression_astc_hdr'

pub type PhysicalDeviceTextureCompressionASTCHDRFeaturesEXT = C.VkPhysicalDeviceTextureCompressionASTCHDRFeatures

pub const ext_astc_decode_mode_spec_version = 1
pub const ext_astc_decode_mode_extension_name = c'VK_EXT_astc_decode_mode'
// ImageViewASTCDecodeModeEXT extends VkImageViewCreateInfo
pub type ImageViewASTCDecodeModeEXT = C.VkImageViewASTCDecodeModeEXT

@[typedef]
pub struct C.VkImageViewASTCDecodeModeEXT {
pub mut:
	sType      StructureType = StructureType.image_view_astc_decode_mode_ext
	pNext      voidptr       = unsafe { nil }
	decodeMode Format
}

// PhysicalDeviceASTCDecodeFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceASTCDecodeFeaturesEXT = C.VkPhysicalDeviceASTCDecodeFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceASTCDecodeFeaturesEXT {
pub mut:
	sType                    StructureType = StructureType.physical_device_astc_decode_features_ext
	pNext                    voidptr       = unsafe { nil }
	decodeModeSharedExponent Bool32
}

pub const ext_pipeline_robustness_spec_version = 1
pub const ext_pipeline_robustness_extension_name = c'VK_EXT_pipeline_robustness'

pub type PipelineRobustnessBufferBehaviorEXT = PipelineRobustnessBufferBehavior

pub type PipelineRobustnessImageBehaviorEXT = PipelineRobustnessImageBehavior

pub type PhysicalDevicePipelineRobustnessFeaturesEXT = C.VkPhysicalDevicePipelineRobustnessFeatures

pub type PhysicalDevicePipelineRobustnessPropertiesEXT = C.VkPhysicalDevicePipelineRobustnessProperties

pub type PipelineRobustnessCreateInfoEXT = C.VkPipelineRobustnessCreateInfo

pub const ext_conditional_rendering_spec_version = 2
pub const ext_conditional_rendering_extension_name = c'VK_EXT_conditional_rendering'

pub enum ConditionalRenderingFlagBitsEXT as u32 {
	inverted     = u32(0x00000001)
	max_enum_ext = max_int
}
pub type ConditionalRenderingFlagsEXT = u32
pub type ConditionalRenderingBeginInfoEXT = C.VkConditionalRenderingBeginInfoEXT

@[typedef]
pub struct C.VkConditionalRenderingBeginInfoEXT {
pub mut:
	sType  StructureType = StructureType.conditional_rendering_begin_info_ext
	pNext  voidptr       = unsafe { nil }
	buffer Buffer
	offset DeviceSize
	flags  ConditionalRenderingFlagsEXT
}

// PhysicalDeviceConditionalRenderingFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceConditionalRenderingFeaturesEXT = C.VkPhysicalDeviceConditionalRenderingFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceConditionalRenderingFeaturesEXT {
pub mut:
	sType                         StructureType = StructureType.physical_device_conditional_rendering_features_ext
	pNext                         voidptr       = unsafe { nil }
	conditionalRendering          Bool32
	inheritedConditionalRendering Bool32
}

// CommandBufferInheritanceConditionalRenderingInfoEXT extends VkCommandBufferInheritanceInfo
pub type CommandBufferInheritanceConditionalRenderingInfoEXT = C.VkCommandBufferInheritanceConditionalRenderingInfoEXT

@[typedef]
pub struct C.VkCommandBufferInheritanceConditionalRenderingInfoEXT {
pub mut:
	sType                      StructureType = StructureType.command_buffer_inheritance_conditional_rendering_info_ext
	pNext                      voidptr       = unsafe { nil }
	conditionalRenderingEnable Bool32
}

@[keep_args_alive]
fn C.vkCmdBeginConditionalRenderingEXT(command_buffer CommandBuffer, p_conditional_rendering_begin &ConditionalRenderingBeginInfoEXT)

pub type PFN_vkCmdBeginConditionalRenderingEXT = fn (command_buffer CommandBuffer, p_conditional_rendering_begin &ConditionalRenderingBeginInfoEXT)

@[inline]
pub fn cmd_begin_conditional_rendering_ext(command_buffer CommandBuffer,
	p_conditional_rendering_begin &ConditionalRenderingBeginInfoEXT) {
	C.vkCmdBeginConditionalRenderingEXT(command_buffer, p_conditional_rendering_begin)
}

@[keep_args_alive]
fn C.vkCmdEndConditionalRenderingEXT(command_buffer CommandBuffer)

pub type PFN_vkCmdEndConditionalRenderingEXT = fn (command_buffer CommandBuffer)

@[inline]
pub fn cmd_end_conditional_rendering_ext(command_buffer CommandBuffer) {
	C.vkCmdEndConditionalRenderingEXT(command_buffer)
}

pub const nv_clip_space_w_scaling_spec_version = 1
pub const nv_clip_space_w_scaling_extension_name = c'VK_NV_clip_space_w_scaling'

pub type ViewportWScalingNV = C.VkViewportWScalingNV

@[typedef]
pub struct C.VkViewportWScalingNV {
pub mut:
	xcoeff f32
	ycoeff f32
}

// PipelineViewportWScalingStateCreateInfoNV extends VkPipelineViewportStateCreateInfo
pub type PipelineViewportWScalingStateCreateInfoNV = C.VkPipelineViewportWScalingStateCreateInfoNV

@[typedef]
pub struct C.VkPipelineViewportWScalingStateCreateInfoNV {
pub mut:
	sType                  StructureType = StructureType.pipeline_viewport_w_scaling_state_create_info_nv
	pNext                  voidptr       = unsafe { nil }
	viewportWScalingEnable Bool32
	viewportCount          u32
	pViewportWScalings     &ViewportWScalingNV
}

@[keep_args_alive]
fn C.vkCmdSetViewportWScalingNV(command_buffer CommandBuffer, first_viewport u32, viewport_count u32, p_viewport_w_scalings &ViewportWScalingNV)

pub type PFN_vkCmdSetViewportWScalingNV = fn (command_buffer CommandBuffer, first_viewport u32, viewport_count u32, p_viewport_w_scalings &ViewportWScalingNV)

@[inline]
pub fn cmd_set_viewport_w_scaling_nv(command_buffer CommandBuffer,
	first_viewport u32,
	viewport_count u32,
	p_viewport_w_scalings &ViewportWScalingNV) {
	C.vkCmdSetViewportWScalingNV(command_buffer, first_viewport, viewport_count, p_viewport_w_scalings)
}

pub const ext_direct_mode_display_spec_version = 1
pub const ext_direct_mode_display_extension_name = c'VK_EXT_direct_mode_display'

@[keep_args_alive]
fn C.vkReleaseDisplayEXT(physical_device PhysicalDevice, display DisplayKHR) Result

pub type PFN_vkReleaseDisplayEXT = fn (physical_device PhysicalDevice, display DisplayKHR) Result

@[inline]
pub fn release_display_ext(physical_device PhysicalDevice,
	display DisplayKHR) Result {
	return C.vkReleaseDisplayEXT(physical_device, display)
}

pub const ext_display_surface_counter_spec_version = 1
pub const ext_display_surface_counter_extension_name = c'VK_EXT_display_surface_counter'

pub enum SurfaceCounterFlagBitsEXT as u32 {
	vblank       = u32(0x00000001)
	max_enum_ext = max_int
}
pub type SurfaceCounterFlagsEXT = u32
pub type SurfaceCapabilities2EXT = C.VkSurfaceCapabilities2EXT

@[typedef]
pub struct C.VkSurfaceCapabilities2EXT {
pub mut:
	sType                    StructureType = StructureType.surface_capabilities2_ext
	pNext                    voidptr       = unsafe { nil }
	minImageCount            u32
	maxImageCount            u32
	currentExtent            Extent2D
	minImageExtent           Extent2D
	maxImageExtent           Extent2D
	maxImageArrayLayers      u32
	supportedTransforms      SurfaceTransformFlagsKHR
	currentTransform         SurfaceTransformFlagBitsKHR
	supportedCompositeAlpha  CompositeAlphaFlagsKHR
	supportedUsageFlags      ImageUsageFlags
	supportedSurfaceCounters SurfaceCounterFlagsEXT
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceSurfaceCapabilities2EXT(physical_device PhysicalDevice, surface SurfaceKHR, mut p_surface_capabilities SurfaceCapabilities2EXT) Result

pub type PFN_vkGetPhysicalDeviceSurfaceCapabilities2EXT = fn (physical_device PhysicalDevice, surface SurfaceKHR, mut p_surface_capabilities SurfaceCapabilities2EXT) Result

@[inline]
pub fn get_physical_device_surface_capabilities2_ext(physical_device PhysicalDevice,
	surface SurfaceKHR,
	mut p_surface_capabilities SurfaceCapabilities2EXT) Result {
	return C.vkGetPhysicalDeviceSurfaceCapabilities2EXT(physical_device, surface, mut
		p_surface_capabilities)
}

pub const ext_display_control_spec_version = 1
pub const ext_display_control_extension_name = c'VK_EXT_display_control'

pub enum DisplayPowerStateEXT as u32 {
	off          = 0
	suspend      = 1
	on           = 2
	max_enum_ext = max_int
}

pub enum DeviceEventTypeEXT as u32 {
	display_hotplug = 0
	max_enum_ext    = max_int
}

pub enum DisplayEventTypeEXT as u32 {
	first_pixel_out = 0
	max_enum_ext    = max_int
}
pub type DisplayPowerInfoEXT = C.VkDisplayPowerInfoEXT

@[typedef]
pub struct C.VkDisplayPowerInfoEXT {
pub mut:
	sType      StructureType = StructureType.display_power_info_ext
	pNext      voidptr       = unsafe { nil }
	powerState DisplayPowerStateEXT
}

pub type DeviceEventInfoEXT = C.VkDeviceEventInfoEXT

@[typedef]
pub struct C.VkDeviceEventInfoEXT {
pub mut:
	sType       StructureType = StructureType.device_event_info_ext
	pNext       voidptr       = unsafe { nil }
	deviceEvent DeviceEventTypeEXT
}

pub type DisplayEventInfoEXT = C.VkDisplayEventInfoEXT

@[typedef]
pub struct C.VkDisplayEventInfoEXT {
pub mut:
	sType        StructureType = StructureType.display_event_info_ext
	pNext        voidptr       = unsafe { nil }
	displayEvent DisplayEventTypeEXT
}

// SwapchainCounterCreateInfoEXT extends VkSwapchainCreateInfoKHR
pub type SwapchainCounterCreateInfoEXT = C.VkSwapchainCounterCreateInfoEXT

@[typedef]
pub struct C.VkSwapchainCounterCreateInfoEXT {
pub mut:
	sType           StructureType = StructureType.swapchain_counter_create_info_ext
	pNext           voidptr       = unsafe { nil }
	surfaceCounters SurfaceCounterFlagsEXT
}

@[keep_args_alive]
fn C.vkDisplayPowerControlEXT(device Device, display DisplayKHR, p_display_power_info &DisplayPowerInfoEXT) Result

pub type PFN_vkDisplayPowerControlEXT = fn (device Device, display DisplayKHR, p_display_power_info &DisplayPowerInfoEXT) Result

@[inline]
pub fn display_power_control_ext(device Device,
	display DisplayKHR,
	p_display_power_info &DisplayPowerInfoEXT) Result {
	return C.vkDisplayPowerControlEXT(device, display, p_display_power_info)
}

@[keep_args_alive]
fn C.vkRegisterDeviceEventEXT(device Device, p_device_event_info &DeviceEventInfoEXT, p_allocator &AllocationCallbacks, p_fence &Fence) Result

pub type PFN_vkRegisterDeviceEventEXT = fn (device Device, p_device_event_info &DeviceEventInfoEXT, p_allocator &AllocationCallbacks, p_fence &Fence) Result

@[inline]
pub fn register_device_event_ext(device Device,
	p_device_event_info &DeviceEventInfoEXT,
	p_allocator &AllocationCallbacks,
	p_fence &Fence) Result {
	return C.vkRegisterDeviceEventEXT(device, p_device_event_info, p_allocator, p_fence)
}

@[keep_args_alive]
fn C.vkRegisterDisplayEventEXT(device Device, display DisplayKHR, p_display_event_info &DisplayEventInfoEXT, p_allocator &AllocationCallbacks, p_fence &Fence) Result

pub type PFN_vkRegisterDisplayEventEXT = fn (device Device, display DisplayKHR, p_display_event_info &DisplayEventInfoEXT, p_allocator &AllocationCallbacks, p_fence &Fence) Result

@[inline]
pub fn register_display_event_ext(device Device,
	display DisplayKHR,
	p_display_event_info &DisplayEventInfoEXT,
	p_allocator &AllocationCallbacks,
	p_fence &Fence) Result {
	return C.vkRegisterDisplayEventEXT(device, display, p_display_event_info, p_allocator,
		p_fence)
}

@[keep_args_alive]
fn C.vkGetSwapchainCounterEXT(device Device, swapchain SwapchainKHR, counter SurfaceCounterFlagBitsEXT, p_counter_value &u64) Result

pub type PFN_vkGetSwapchainCounterEXT = fn (device Device, swapchain SwapchainKHR, counter SurfaceCounterFlagBitsEXT, p_counter_value &u64) Result

@[inline]
pub fn get_swapchain_counter_ext(device Device,
	swapchain SwapchainKHR,
	counter SurfaceCounterFlagBitsEXT,
	p_counter_value &u64) Result {
	return C.vkGetSwapchainCounterEXT(device, swapchain, counter, p_counter_value)
}

pub const google_display_timing_spec_version = 1
pub const google_display_timing_extension_name = c'VK_GOOGE_display_timing'

pub type RefreshCycleDurationGOOGLE = C.VkRefreshCycleDurationGOOGLE

@[typedef]
pub struct C.VkRefreshCycleDurationGOOGLE {
pub mut:
	refreshDuration u64
}

pub type PastPresentationTimingGOOGLE = C.VkPastPresentationTimingGOOGLE

@[typedef]
pub struct C.VkPastPresentationTimingGOOGLE {
pub mut:
	presentID           u32
	desiredPresentTime  u64
	actualPresentTime   u64
	earliestPresentTime u64
	presentMargin       u64
}

pub type PresentTimeGOOGLE = C.VkPresentTimeGOOGLE

@[typedef]
pub struct C.VkPresentTimeGOOGLE {
pub mut:
	presentID          u32
	desiredPresentTime u64
}

// PresentTimesInfoGOOGLE extends VkPresentInfoKHR
pub type PresentTimesInfoGOOGLE = C.VkPresentTimesInfoGOOGLE

@[typedef]
pub struct C.VkPresentTimesInfoGOOGLE {
pub mut:
	sType          StructureType = StructureType.present_times_info_google
	pNext          voidptr       = unsafe { nil }
	swapchainCount u32
	pTimes         &PresentTimeGOOGLE
}

@[keep_args_alive]
fn C.vkGetRefreshCycleDurationGOOGLE(device Device, swapchain SwapchainKHR, mut p_display_timing_properties RefreshCycleDurationGOOGLE) Result

pub type PFN_vkGetRefreshCycleDurationGOOGLE = fn (device Device, swapchain SwapchainKHR, mut p_display_timing_properties RefreshCycleDurationGOOGLE) Result

@[inline]
pub fn get_refresh_cycle_duration_google(device Device,
	swapchain SwapchainKHR,
	mut p_display_timing_properties RefreshCycleDurationGOOGLE) Result {
	return C.vkGetRefreshCycleDurationGOOGLE(device, swapchain, mut p_display_timing_properties)
}

@[keep_args_alive]
fn C.vkGetPastPresentationTimingGOOGLE(device Device, swapchain SwapchainKHR, p_presentation_timing_count &u32, mut p_presentation_timings PastPresentationTimingGOOGLE) Result

pub type PFN_vkGetPastPresentationTimingGOOGLE = fn (device Device, swapchain SwapchainKHR, p_presentation_timing_count &u32, mut p_presentation_timings PastPresentationTimingGOOGLE) Result

@[inline]
pub fn get_past_presentation_timing_google(device Device,
	swapchain SwapchainKHR,
	p_presentation_timing_count &u32,
	mut p_presentation_timings PastPresentationTimingGOOGLE) Result {
	return C.vkGetPastPresentationTimingGOOGLE(device, swapchain, p_presentation_timing_count, mut
		p_presentation_timings)
}

pub const nv_sample_mask_override_coverage_spec_version = 1
pub const nv_sample_mask_override_coverage_extension_name = c'VK_NV_sample_mask_override_coverage'

pub const nv_geometry_shader_passthrough_spec_version = 1
pub const nv_geometry_shader_passthrough_extension_name = c'VK_NV_geometry_shader_passthrough'

pub const nv_viewport_array_2_spec_version = 1
pub const nv_viewport_array_2_extension_name = c'VK_NV_viewport_array2'
// VK_NV_VIEWPORT_ARRAY2_SPEC_VERSION is a deprecated alias
pub const nv_viewport_array2_spec_version = nv_viewport_array_2_spec_version
// VK_NV_VIEWPORT_ARRAY2_EXTENSION_NAME is a deprecated alias
pub const nv_viewport_array2_extension_name = nv_viewport_array_2_extension_name

pub const nvx_multiview_per_view_attributes_spec_version = 1
pub const nvx_multiview_per_view_attributes_extension_name = c'VK_NVX_multiview_per_view_attributes'
// PhysicalDeviceMultiviewPerViewAttributesPropertiesNVX extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMultiviewPerViewAttributesPropertiesNVX = C.VkPhysicalDeviceMultiviewPerViewAttributesPropertiesNVX

@[typedef]
pub struct C.VkPhysicalDeviceMultiviewPerViewAttributesPropertiesNVX {
pub mut:
	sType                        StructureType = StructureType.physical_device_multiview_per_view_attributes_properties_nvx
	pNext                        voidptr       = unsafe { nil }
	perViewPositionAllComponents Bool32
}

// MultiviewPerViewAttributesInfoNVX extends VkCommandBufferInheritanceInfo,VkGraphicsPipelineCreateInfo,VkRenderingInfo
pub type MultiviewPerViewAttributesInfoNVX = C.VkMultiviewPerViewAttributesInfoNVX

@[typedef]
pub struct C.VkMultiviewPerViewAttributesInfoNVX {
pub mut:
	sType                          StructureType = StructureType.multiview_per_view_attributes_info_nvx
	pNext                          voidptr       = unsafe { nil }
	perViewAttributes              Bool32
	perViewAttributesPositionXOnly Bool32
}

pub const nv_viewport_swizzle_spec_version = 1
pub const nv_viewport_swizzle_extension_name = c'VK_NV_viewport_swizzle'

pub enum ViewportCoordinateSwizzleNV as u32 {
	positive_x  = 0
	negative_x  = 1
	positive_y  = 2
	negative_y  = 3
	positive_z  = 4
	negative_z  = 5
	positive_w  = 6
	negative_w  = 7
	max_enum_nv = max_int
}
pub type PipelineViewportSwizzleStateCreateFlagsNV = u32
pub type ViewportSwizzleNV = C.VkViewportSwizzleNV

@[typedef]
pub struct C.VkViewportSwizzleNV {
pub mut:
	x ViewportCoordinateSwizzleNV
	y ViewportCoordinateSwizzleNV
	z ViewportCoordinateSwizzleNV
	w ViewportCoordinateSwizzleNV
}

// PipelineViewportSwizzleStateCreateInfoNV extends VkPipelineViewportStateCreateInfo
pub type PipelineViewportSwizzleStateCreateInfoNV = C.VkPipelineViewportSwizzleStateCreateInfoNV

@[typedef]
pub struct C.VkPipelineViewportSwizzleStateCreateInfoNV {
pub mut:
	sType             StructureType = StructureType.pipeline_viewport_swizzle_state_create_info_nv
	pNext             voidptr       = unsafe { nil }
	flags             PipelineViewportSwizzleStateCreateFlagsNV
	viewportCount     u32
	pViewportSwizzles &ViewportSwizzleNV
}

pub const ext_discard_rectangles_spec_version = 2
pub const ext_discard_rectangles_extension_name = c'VK_EXT_discard_rectangles'

pub enum DiscardRectangleModeEXT as u32 {
	inclusive    = 0
	exclusive    = 1
	max_enum_ext = max_int
}
pub type PipelineDiscardRectangleStateCreateFlagsEXT = u32

// PhysicalDeviceDiscardRectanglePropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceDiscardRectanglePropertiesEXT = C.VkPhysicalDeviceDiscardRectanglePropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDiscardRectanglePropertiesEXT {
pub mut:
	sType                StructureType = StructureType.physical_device_discard_rectangle_properties_ext
	pNext                voidptr       = unsafe { nil }
	maxDiscardRectangles u32
}

// PipelineDiscardRectangleStateCreateInfoEXT extends VkGraphicsPipelineCreateInfo
pub type PipelineDiscardRectangleStateCreateInfoEXT = C.VkPipelineDiscardRectangleStateCreateInfoEXT

@[typedef]
pub struct C.VkPipelineDiscardRectangleStateCreateInfoEXT {
pub mut:
	sType                 StructureType = StructureType.pipeline_discard_rectangle_state_create_info_ext
	pNext                 voidptr       = unsafe { nil }
	flags                 PipelineDiscardRectangleStateCreateFlagsEXT
	discardRectangleMode  DiscardRectangleModeEXT
	discardRectangleCount u32
	pDiscardRectangles    &Rect2D
}

@[keep_args_alive]
fn C.vkCmdSetDiscardRectangleEXT(command_buffer CommandBuffer, first_discard_rectangle u32, discard_rectangle_count u32, p_discard_rectangles &Rect2D)

pub type PFN_vkCmdSetDiscardRectangleEXT = fn (command_buffer CommandBuffer, first_discard_rectangle u32, discard_rectangle_count u32, p_discard_rectangles &Rect2D)

@[inline]
pub fn cmd_set_discard_rectangle_ext(command_buffer CommandBuffer,
	first_discard_rectangle u32,
	discard_rectangle_count u32,
	p_discard_rectangles &Rect2D) {
	C.vkCmdSetDiscardRectangleEXT(command_buffer, first_discard_rectangle, discard_rectangle_count,
		p_discard_rectangles)
}

@[keep_args_alive]
fn C.vkCmdSetDiscardRectangleEnableEXT(command_buffer CommandBuffer, discard_rectangle_enable Bool32)

pub type PFN_vkCmdSetDiscardRectangleEnableEXT = fn (command_buffer CommandBuffer, discard_rectangle_enable Bool32)

@[inline]
pub fn cmd_set_discard_rectangle_enable_ext(command_buffer CommandBuffer,
	discard_rectangle_enable Bool32) {
	C.vkCmdSetDiscardRectangleEnableEXT(command_buffer, discard_rectangle_enable)
}

@[keep_args_alive]
fn C.vkCmdSetDiscardRectangleModeEXT(command_buffer CommandBuffer, discard_rectangle_mode DiscardRectangleModeEXT)

pub type PFN_vkCmdSetDiscardRectangleModeEXT = fn (command_buffer CommandBuffer, discard_rectangle_mode DiscardRectangleModeEXT)

@[inline]
pub fn cmd_set_discard_rectangle_mode_ext(command_buffer CommandBuffer,
	discard_rectangle_mode DiscardRectangleModeEXT) {
	C.vkCmdSetDiscardRectangleModeEXT(command_buffer, discard_rectangle_mode)
}

pub const ext_conservative_rasterization_spec_version = 1
pub const ext_conservative_rasterization_extension_name = c'VK_EXT_conservative_rasterization'

pub enum ConservativeRasterizationModeEXT as u32 {
	disabled      = 0
	overestimate  = 1
	underestimate = 2
	max_enum_ext  = max_int
}
pub type PipelineRasterizationConservativeStateCreateFlagsEXT = u32

// PhysicalDeviceConservativeRasterizationPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceConservativeRasterizationPropertiesEXT = C.VkPhysicalDeviceConservativeRasterizationPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceConservativeRasterizationPropertiesEXT {
pub mut:
	sType                                       StructureType = StructureType.physical_device_conservative_rasterization_properties_ext
	pNext                                       voidptr       = unsafe { nil }
	primitiveOverestimationSize                 f32
	maxExtraPrimitiveOverestimationSize         f32
	extraPrimitiveOverestimationSizeGranularity f32
	primitiveUnderestimation                    Bool32
	conservativePointAndLineRasterization       Bool32
	degenerateTrianglesRasterized               Bool32
	degenerateLinesRasterized                   Bool32
	fullyCoveredFragmentShaderInputVariable     Bool32
	conservativeRasterizationPostDepthCoverage  Bool32
}

// PipelineRasterizationConservativeStateCreateInfoEXT extends VkPipelineRasterizationStateCreateInfo
pub type PipelineRasterizationConservativeStateCreateInfoEXT = C.VkPipelineRasterizationConservativeStateCreateInfoEXT

@[typedef]
pub struct C.VkPipelineRasterizationConservativeStateCreateInfoEXT {
pub mut:
	sType                            StructureType = StructureType.pipeline_rasterization_conservative_state_create_info_ext
	pNext                            voidptr       = unsafe { nil }
	flags                            PipelineRasterizationConservativeStateCreateFlagsEXT
	conservativeRasterizationMode    ConservativeRasterizationModeEXT
	extraPrimitiveOverestimationSize f32
}

pub const ext_depth_clip_enable_spec_version = 1
pub const ext_depth_clip_enable_extension_name = c'VK_EXT_depth_clip_enable'

pub type PipelineRasterizationDepthClipStateCreateFlagsEXT = u32

// PhysicalDeviceDepthClipEnableFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDepthClipEnableFeaturesEXT = C.VkPhysicalDeviceDepthClipEnableFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDepthClipEnableFeaturesEXT {
pub mut:
	sType           StructureType = StructureType.physical_device_depth_clip_enable_features_ext
	pNext           voidptr       = unsafe { nil }
	depthClipEnable Bool32
}

// PipelineRasterizationDepthClipStateCreateInfoEXT extends VkPipelineRasterizationStateCreateInfo
pub type PipelineRasterizationDepthClipStateCreateInfoEXT = C.VkPipelineRasterizationDepthClipStateCreateInfoEXT

@[typedef]
pub struct C.VkPipelineRasterizationDepthClipStateCreateInfoEXT {
pub mut:
	sType           StructureType = StructureType.pipeline_rasterization_depth_clip_state_create_info_ext
	pNext           voidptr       = unsafe { nil }
	flags           PipelineRasterizationDepthClipStateCreateFlagsEXT
	depthClipEnable Bool32
}

pub const ext_swapchain_color_space_spec_version = 5
pub const ext_swapchain_color_space_extension_name = c'VK_EXT_swapchain_colorspace'

pub const ext_hdr_metadata_spec_version = 3
pub const ext_hdr_metadata_extension_name = c'VK_EXT_hdr_metadata'

pub type XYColorEXT = C.VkXYColorEXT

@[typedef]
pub struct C.VkXYColorEXT {
pub mut:
	x f32
	y f32
}

pub type HdrMetadataEXT = C.VkHdrMetadataEXT

@[typedef]
pub struct C.VkHdrMetadataEXT {
pub mut:
	sType                     StructureType = StructureType.hdr_metadata_ext
	pNext                     voidptr       = unsafe { nil }
	displayPrimaryRed         XYColorEXT
	displayPrimaryGreen       XYColorEXT
	displayPrimaryBlue        XYColorEXT
	whitePoint                XYColorEXT
	maxLuminance              f32
	minLuminance              f32
	maxContentLightLevel      f32
	maxFrameAverageLightLevel f32
}

@[keep_args_alive]
fn C.vkSetHdrMetadataEXT(device Device, swapchain_count u32, p_swapchains &SwapchainKHR, p_metadata &HdrMetadataEXT)

pub type PFN_vkSetHdrMetadataEXT = fn (device Device, swapchain_count u32, p_swapchains &SwapchainKHR, p_metadata &HdrMetadataEXT)

@[inline]
pub fn set_hdr_metadata_ext(device Device,
	swapchain_count u32,
	p_swapchains &SwapchainKHR,
	p_metadata &HdrMetadataEXT) {
	C.vkSetHdrMetadataEXT(device, swapchain_count, p_swapchains, p_metadata)
}

pub const img_relaxed_line_rasterization_spec_version = 1
pub const img_relaxed_line_rasterization_extension_name = c'VK_IMG_relaxed_line_rasterization'
// PhysicalDeviceRelaxedLineRasterizationFeaturesIMG extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRelaxedLineRasterizationFeaturesIMG = C.VkPhysicalDeviceRelaxedLineRasterizationFeaturesIMG

@[typedef]
pub struct C.VkPhysicalDeviceRelaxedLineRasterizationFeaturesIMG {
pub mut:
	sType                    StructureType = StructureType.physical_device_relaxed_line_rasterization_features_img
	pNext                    voidptr       = unsafe { nil }
	relaxedLineRasterization Bool32
}

pub const ext_external_memory_dma_buf_spec_version = 1
pub const ext_external_memory_dma_buf_extension_name = c'VK_EXT_external_memory_dma_buf'

pub const ext_queue_family_foreign_spec_version = 1
pub const ext_queue_family_foreign_extension_name = c'VK_EXT_queue_family_foreign'
pub const queue_family_foreign_ext = ~u32(2)

// Pointer to VkDebugUtilsMessengerEXT_T
pub type DebugUtilsMessengerEXT = voidptr

pub const ext_debug_utils_spec_version = 2
pub const ext_debug_utils_extension_name = c'VK_EXT_debug_utils'

pub type DebugUtilsMessengerCallbackDataFlagsEXT = u32

pub enum DebugUtilsMessageSeverityFlagBitsEXT as u32 {
	verbose      = u32(0x00000001)
	info         = u32(0x00000010)
	warning      = u32(0x00000100)
	error        = u32(0x00001000)
	max_enum_ext = max_int
}

pub enum DebugUtilsMessageTypeFlagBitsEXT as u32 {
	general                = u32(0x00000001)
	validation             = u32(0x00000002)
	performance            = u32(0x00000004)
	device_address_binding = u32(0x00000008)
	max_enum_ext           = max_int
}
pub type DebugUtilsMessageTypeFlagsEXT = u32
pub type DebugUtilsMessageSeverityFlagsEXT = u32
pub type DebugUtilsMessengerCreateFlagsEXT = u32
pub type DebugUtilsLabelEXT = C.VkDebugUtilsLabelEXT

@[typedef]
pub struct C.VkDebugUtilsLabelEXT {
pub mut:
	sType      StructureType = StructureType.debug_utils_label_ext
	pNext      voidptr       = unsafe { nil }
	pLabelName &char
	color      [4]f32
}

// DebugUtilsObjectNameInfoEXT extends VkPipelineShaderStageCreateInfo
pub type DebugUtilsObjectNameInfoEXT = C.VkDebugUtilsObjectNameInfoEXT

@[typedef]
pub struct C.VkDebugUtilsObjectNameInfoEXT {
pub mut:
	sType        StructureType = StructureType.debug_utils_object_name_info_ext
	pNext        voidptr       = unsafe { nil }
	objectType   ObjectType
	objectHandle u64
	pObjectName  &char
}

pub type DebugUtilsMessengerCallbackDataEXT = C.VkDebugUtilsMessengerCallbackDataEXT

@[typedef]
pub struct C.VkDebugUtilsMessengerCallbackDataEXT {
pub mut:
	sType            StructureType = StructureType.debug_utils_messenger_callback_data_ext
	pNext            voidptr       = unsafe { nil }
	flags            DebugUtilsMessengerCallbackDataFlagsEXT
	pMessageIdName   &char
	messageIdNumber  i32
	pMessage         &char
	queueLabelCount  u32
	pQueueLabels     &DebugUtilsLabelEXT
	cmdBufLabelCount u32
	pCmdBufLabels    &DebugUtilsLabelEXT
	objectCount      u32
	pObjects         &DebugUtilsObjectNameInfoEXT
}

pub type PFN_vkDebugUtilsMessengerCallbackEXT = fn (DebugUtilsMessageSeverityFlagBitsEXT, DebugUtilsMessageTypeFlagsEXT, &DebugUtilsMessengerCallbackDataEXT, voidptr)

// DebugUtilsMessengerCreateInfoEXT extends VkInstanceCreateInfo
pub type DebugUtilsMessengerCreateInfoEXT = C.VkDebugUtilsMessengerCreateInfoEXT

@[typedef]
pub struct C.VkDebugUtilsMessengerCreateInfoEXT {
pub mut:
	sType           StructureType = StructureType.debug_utils_messenger_create_info_ext
	pNext           voidptr       = unsafe { nil }
	flags           DebugUtilsMessengerCreateFlagsEXT
	messageSeverity DebugUtilsMessageSeverityFlagsEXT
	messageType     DebugUtilsMessageTypeFlagsEXT
	pfnUserCallback PFN_vkDebugUtilsMessengerCallbackEXT = unsafe { nil }
	pUserData       voidptr = unsafe { nil }
}

pub type DebugUtilsObjectTagInfoEXT = C.VkDebugUtilsObjectTagInfoEXT

@[typedef]
pub struct C.VkDebugUtilsObjectTagInfoEXT {
pub mut:
	sType        StructureType = StructureType.debug_utils_object_tag_info_ext
	pNext        voidptr       = unsafe { nil }
	objectType   ObjectType
	objectHandle u64
	tagName      u64
	tagSize      usize
	pTag         voidptr
}

@[keep_args_alive]
fn C.vkSetDebugUtilsObjectNameEXT(device Device, p_name_info &DebugUtilsObjectNameInfoEXT) Result

pub type PFN_vkSetDebugUtilsObjectNameEXT = fn (device Device, p_name_info &DebugUtilsObjectNameInfoEXT) Result

@[inline]
pub fn set_debug_utils_object_name_ext(device Device,
	p_name_info &DebugUtilsObjectNameInfoEXT) Result {
	return C.vkSetDebugUtilsObjectNameEXT(device, p_name_info)
}

@[keep_args_alive]
fn C.vkSetDebugUtilsObjectTagEXT(device Device, p_tag_info &DebugUtilsObjectTagInfoEXT) Result

pub type PFN_vkSetDebugUtilsObjectTagEXT = fn (device Device, p_tag_info &DebugUtilsObjectTagInfoEXT) Result

@[inline]
pub fn set_debug_utils_object_tag_ext(device Device,
	p_tag_info &DebugUtilsObjectTagInfoEXT) Result {
	return C.vkSetDebugUtilsObjectTagEXT(device, p_tag_info)
}

@[keep_args_alive]
fn C.vkQueueBeginDebugUtilsLabelEXT(queue Queue, p_label_info &DebugUtilsLabelEXT)

pub type PFN_vkQueueBeginDebugUtilsLabelEXT = fn (queue Queue, p_label_info &DebugUtilsLabelEXT)

@[inline]
pub fn queue_begin_debug_utils_label_ext(queue Queue,
	p_label_info &DebugUtilsLabelEXT) {
	C.vkQueueBeginDebugUtilsLabelEXT(queue, p_label_info)
}

@[keep_args_alive]
fn C.vkQueueEndDebugUtilsLabelEXT(queue Queue)

pub type PFN_vkQueueEndDebugUtilsLabelEXT = fn (queue Queue)

@[inline]
pub fn queue_end_debug_utils_label_ext(queue Queue) {
	C.vkQueueEndDebugUtilsLabelEXT(queue)
}

@[keep_args_alive]
fn C.vkQueueInsertDebugUtilsLabelEXT(queue Queue, p_label_info &DebugUtilsLabelEXT)

pub type PFN_vkQueueInsertDebugUtilsLabelEXT = fn (queue Queue, p_label_info &DebugUtilsLabelEXT)

@[inline]
pub fn queue_insert_debug_utils_label_ext(queue Queue,
	p_label_info &DebugUtilsLabelEXT) {
	C.vkQueueInsertDebugUtilsLabelEXT(queue, p_label_info)
}

@[keep_args_alive]
fn C.vkCmdBeginDebugUtilsLabelEXT(command_buffer CommandBuffer, p_label_info &DebugUtilsLabelEXT)

pub type PFN_vkCmdBeginDebugUtilsLabelEXT = fn (command_buffer CommandBuffer, p_label_info &DebugUtilsLabelEXT)

@[inline]
pub fn cmd_begin_debug_utils_label_ext(command_buffer CommandBuffer,
	p_label_info &DebugUtilsLabelEXT) {
	C.vkCmdBeginDebugUtilsLabelEXT(command_buffer, p_label_info)
}

@[keep_args_alive]
fn C.vkCmdEndDebugUtilsLabelEXT(command_buffer CommandBuffer)

pub type PFN_vkCmdEndDebugUtilsLabelEXT = fn (command_buffer CommandBuffer)

@[inline]
pub fn cmd_end_debug_utils_label_ext(command_buffer CommandBuffer) {
	C.vkCmdEndDebugUtilsLabelEXT(command_buffer)
}

@[keep_args_alive]
fn C.vkCmdInsertDebugUtilsLabelEXT(command_buffer CommandBuffer, p_label_info &DebugUtilsLabelEXT)

pub type PFN_vkCmdInsertDebugUtilsLabelEXT = fn (command_buffer CommandBuffer, p_label_info &DebugUtilsLabelEXT)

@[inline]
pub fn cmd_insert_debug_utils_label_ext(command_buffer CommandBuffer,
	p_label_info &DebugUtilsLabelEXT) {
	C.vkCmdInsertDebugUtilsLabelEXT(command_buffer, p_label_info)
}

@[keep_args_alive]
fn C.vkCreateDebugUtilsMessengerEXT(instance Instance, p_create_info &DebugUtilsMessengerCreateInfoEXT, p_allocator &AllocationCallbacks, p_messenger &DebugUtilsMessengerEXT) Result

pub type PFN_vkCreateDebugUtilsMessengerEXT = fn (instance Instance, p_create_info &DebugUtilsMessengerCreateInfoEXT, p_allocator &AllocationCallbacks, p_messenger &DebugUtilsMessengerEXT) Result

@[inline]
pub fn create_debug_utils_messenger_ext(instance Instance,
	p_create_info &DebugUtilsMessengerCreateInfoEXT,
	p_allocator &AllocationCallbacks,
	p_messenger &DebugUtilsMessengerEXT) Result {
	return C.vkCreateDebugUtilsMessengerEXT(instance, p_create_info, p_allocator, p_messenger)
}

@[keep_args_alive]
fn C.vkDestroyDebugUtilsMessengerEXT(instance Instance, messenger DebugUtilsMessengerEXT, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyDebugUtilsMessengerEXT = fn (instance Instance, messenger DebugUtilsMessengerEXT, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_debug_utils_messenger_ext(instance Instance,
	messenger DebugUtilsMessengerEXT,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyDebugUtilsMessengerEXT(instance, messenger, p_allocator)
}

@[keep_args_alive]
fn C.vkSubmitDebugUtilsMessageEXT(instance Instance, message_severity DebugUtilsMessageSeverityFlagBitsEXT, message_types DebugUtilsMessageTypeFlagsEXT, p_callback_data &DebugUtilsMessengerCallbackDataEXT)

pub type PFN_vkSubmitDebugUtilsMessageEXT = fn (instance Instance, message_severity DebugUtilsMessageSeverityFlagBitsEXT, message_types DebugUtilsMessageTypeFlagsEXT, p_callback_data &DebugUtilsMessengerCallbackDataEXT)

@[inline]
pub fn submit_debug_utils_message_ext(instance Instance,
	message_severity DebugUtilsMessageSeverityFlagBitsEXT,
	message_types DebugUtilsMessageTypeFlagsEXT,
	p_callback_data &DebugUtilsMessengerCallbackDataEXT) {
	C.vkSubmitDebugUtilsMessageEXT(instance, message_severity, message_types, p_callback_data)
}

pub const ext_sampler_filter_minmax_spec_version = 2
pub const ext_sampler_filter_minmax_extension_name = c'VK_EXT_sampler_filter_minmax'

pub type SamplerReductionModeEXT = SamplerReductionMode

pub type SamplerReductionModeCreateInfoEXT = C.VkSamplerReductionModeCreateInfo

pub type PhysicalDeviceSamplerFilterMinmaxPropertiesEXT = C.VkPhysicalDeviceSamplerFilterMinmaxProperties

pub const amd_gpu_shader_int16_spec_version = 2
pub const amd_gpu_shader_int16_extension_name = c'VK_AMD_gpu_shader_int16'

pub const amd_mixed_attachment_samples_spec_version = 1
pub const amd_mixed_attachment_samples_extension_name = c'VK_AMD_mixed_attachment_samples'
// AttachmentSampleCountInfoAMD extends VkCommandBufferInheritanceInfo,VkGraphicsPipelineCreateInfo
pub type AttachmentSampleCountInfoAMD = C.VkAttachmentSampleCountInfoAMD

@[typedef]
pub struct C.VkAttachmentSampleCountInfoAMD {
pub mut:
	sType                         StructureType = StructureType.attachment_sample_count_info_amd
	pNext                         voidptr       = unsafe { nil }
	colorAttachmentCount          u32
	pColorAttachmentSamples       &SampleCountFlagBits
	depthStencilAttachmentSamples SampleCountFlagBits
}

pub const amd_shader_fragment_mask_spec_version = 1
pub const amd_shader_fragment_mask_extension_name = c'VK_AMD_shader_fragment_mask'

pub const ext_inline_uniform_block_spec_version = 1
pub const ext_inline_uniform_block_extension_name = c'VK_EXT_inline_uniform_block'

pub type PhysicalDeviceInlineUniformBlockFeaturesEXT = C.VkPhysicalDeviceInlineUniformBlockFeatures

pub type PhysicalDeviceInlineUniformBlockPropertiesEXT = C.VkPhysicalDeviceInlineUniformBlockProperties

pub type WriteDescriptorSetInlineUniformBlockEXT = C.VkWriteDescriptorSetInlineUniformBlock

pub type DescriptorPoolInlineUniformBlockCreateInfoEXT = C.VkDescriptorPoolInlineUniformBlockCreateInfo

pub const ext_shader_stencil_export_spec_version = 1
pub const ext_shader_stencil_export_extension_name = c'VK_EXT_shader_stencil_export'

pub const ext_sample_locations_spec_version = 1
pub const ext_sample_locations_extension_name = c'VK_EXT_sample_locations'

pub type SampleLocationEXT = C.VkSampleLocationEXT

@[typedef]
pub struct C.VkSampleLocationEXT {
pub mut:
	x f32
	y f32
}

// SampleLocationsInfoEXT extends VkImageMemoryBarrier,VkImageMemoryBarrier2
pub type SampleLocationsInfoEXT = C.VkSampleLocationsInfoEXT

@[typedef]
pub struct C.VkSampleLocationsInfoEXT {
pub mut:
	sType                   StructureType = StructureType.sample_locations_info_ext
	pNext                   voidptr       = unsafe { nil }
	sampleLocationsPerPixel SampleCountFlagBits
	sampleLocationGridSize  Extent2D
	sampleLocationsCount    u32
	pSampleLocations        &SampleLocationEXT
}

pub type AttachmentSampleLocationsEXT = C.VkAttachmentSampleLocationsEXT

@[typedef]
pub struct C.VkAttachmentSampleLocationsEXT {
pub mut:
	attachmentIndex     u32
	sampleLocationsInfo SampleLocationsInfoEXT
}

pub type SubpassSampleLocationsEXT = C.VkSubpassSampleLocationsEXT

@[typedef]
pub struct C.VkSubpassSampleLocationsEXT {
pub mut:
	subpassIndex        u32
	sampleLocationsInfo SampleLocationsInfoEXT
}

// RenderPassSampleLocationsBeginInfoEXT extends VkRenderPassBeginInfo
pub type RenderPassSampleLocationsBeginInfoEXT = C.VkRenderPassSampleLocationsBeginInfoEXT

@[typedef]
pub struct C.VkRenderPassSampleLocationsBeginInfoEXT {
pub mut:
	sType                                 StructureType = StructureType.render_pass_sample_locations_begin_info_ext
	pNext                                 voidptr       = unsafe { nil }
	attachmentInitialSampleLocationsCount u32
	pAttachmentInitialSampleLocations     &AttachmentSampleLocationsEXT
	postSubpassSampleLocationsCount       u32
	pPostSubpassSampleLocations           &SubpassSampleLocationsEXT
}

// PipelineSampleLocationsStateCreateInfoEXT extends VkPipelineMultisampleStateCreateInfo
pub type PipelineSampleLocationsStateCreateInfoEXT = C.VkPipelineSampleLocationsStateCreateInfoEXT

@[typedef]
pub struct C.VkPipelineSampleLocationsStateCreateInfoEXT {
pub mut:
	sType                 StructureType = StructureType.pipeline_sample_locations_state_create_info_ext
	pNext                 voidptr       = unsafe { nil }
	sampleLocationsEnable Bool32
	sampleLocationsInfo   SampleLocationsInfoEXT
}

// PhysicalDeviceSampleLocationsPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceSampleLocationsPropertiesEXT = C.VkPhysicalDeviceSampleLocationsPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceSampleLocationsPropertiesEXT {
pub mut:
	sType                         StructureType = StructureType.physical_device_sample_locations_properties_ext
	pNext                         voidptr       = unsafe { nil }
	sampleLocationSampleCounts    SampleCountFlags
	maxSampleLocationGridSize     Extent2D
	sampleLocationCoordinateRange [2]f32
	sampleLocationSubPixelBits    u32
	variableSampleLocations       Bool32
}

pub type MultisamplePropertiesEXT = C.VkMultisamplePropertiesEXT

@[typedef]
pub struct C.VkMultisamplePropertiesEXT {
pub mut:
	sType                     StructureType = StructureType.multisample_properties_ext
	pNext                     voidptr       = unsafe { nil }
	maxSampleLocationGridSize Extent2D
}

@[keep_args_alive]
fn C.vkCmdSetSampleLocationsEXT(command_buffer CommandBuffer, p_sample_locations_info &SampleLocationsInfoEXT)

pub type PFN_vkCmdSetSampleLocationsEXT = fn (command_buffer CommandBuffer, p_sample_locations_info &SampleLocationsInfoEXT)

@[inline]
pub fn cmd_set_sample_locations_ext(command_buffer CommandBuffer,
	p_sample_locations_info &SampleLocationsInfoEXT) {
	C.vkCmdSetSampleLocationsEXT(command_buffer, p_sample_locations_info)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceMultisamplePropertiesEXT(physical_device PhysicalDevice, samples SampleCountFlagBits, mut p_multisample_properties MultisamplePropertiesEXT)

pub type PFN_vkGetPhysicalDeviceMultisamplePropertiesEXT = fn (physical_device PhysicalDevice, samples SampleCountFlagBits, mut p_multisample_properties MultisamplePropertiesEXT)

@[inline]
pub fn get_physical_device_multisample_properties_ext(physical_device PhysicalDevice,
	samples SampleCountFlagBits,
	mut p_multisample_properties MultisamplePropertiesEXT) {
	C.vkGetPhysicalDeviceMultisamplePropertiesEXT(physical_device, samples, mut p_multisample_properties)
}

pub const ext_blend_operation_advanced_spec_version = 2
pub const ext_blend_operation_advanced_extension_name = c'VK_EXT_blend_operation_advanced'

pub enum BlendOverlapEXT as u32 {
	uncorrelated = 0
	disjoint     = 1
	conjoint     = 2
	max_enum_ext = max_int
}
// PhysicalDeviceBlendOperationAdvancedFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceBlendOperationAdvancedFeaturesEXT = C.VkPhysicalDeviceBlendOperationAdvancedFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceBlendOperationAdvancedFeaturesEXT {
pub mut:
	sType                           StructureType = StructureType.physical_device_blend_operation_advanced_features_ext
	pNext                           voidptr       = unsafe { nil }
	advancedBlendCoherentOperations Bool32
}

// PhysicalDeviceBlendOperationAdvancedPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceBlendOperationAdvancedPropertiesEXT = C.VkPhysicalDeviceBlendOperationAdvancedPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceBlendOperationAdvancedPropertiesEXT {
pub mut:
	sType                                 StructureType = StructureType.physical_device_blend_operation_advanced_properties_ext
	pNext                                 voidptr       = unsafe { nil }
	advancedBlendMaxColorAttachments      u32
	advancedBlendIndependentBlend         Bool32
	advancedBlendNonPremultipliedSrcColor Bool32
	advancedBlendNonPremultipliedDstColor Bool32
	advancedBlendCorrelatedOverlap        Bool32
	advancedBlendAllOperations            Bool32
}

// PipelineColorBlendAdvancedStateCreateInfoEXT extends VkPipelineColorBlendStateCreateInfo
pub type PipelineColorBlendAdvancedStateCreateInfoEXT = C.VkPipelineColorBlendAdvancedStateCreateInfoEXT

@[typedef]
pub struct C.VkPipelineColorBlendAdvancedStateCreateInfoEXT {
pub mut:
	sType            StructureType = StructureType.pipeline_color_blend_advanced_state_create_info_ext
	pNext            voidptr       = unsafe { nil }
	srcPremultiplied Bool32
	dstPremultiplied Bool32
	blendOverlap     BlendOverlapEXT
}

pub const nv_fragment_coverage_to_color_spec_version = 1
pub const nv_fragment_coverage_to_color_extension_name = c'VK_NV_fragment_coverage_to_color'

pub type PipelineCoverageToColorStateCreateFlagsNV = u32

// PipelineCoverageToColorStateCreateInfoNV extends VkPipelineMultisampleStateCreateInfo
pub type PipelineCoverageToColorStateCreateInfoNV = C.VkPipelineCoverageToColorStateCreateInfoNV

@[typedef]
pub struct C.VkPipelineCoverageToColorStateCreateInfoNV {
pub mut:
	sType                   StructureType = StructureType.pipeline_coverage_to_color_state_create_info_nv
	pNext                   voidptr       = unsafe { nil }
	flags                   PipelineCoverageToColorStateCreateFlagsNV
	coverageToColorEnable   Bool32
	coverageToColorLocation u32
}

pub const nv_framebuffer_mixed_samples_spec_version = 1
pub const nv_framebuffer_mixed_samples_extension_name = c'VK_NV_framebuffer_mixed_samples'

pub enum CoverageModulationModeNV as u32 {
	none        = 0
	rgb         = 1
	alpha       = 2
	rgba        = 3
	max_enum_nv = max_int
}
pub type PipelineCoverageModulationStateCreateFlagsNV = u32

// PipelineCoverageModulationStateCreateInfoNV extends VkPipelineMultisampleStateCreateInfo
pub type PipelineCoverageModulationStateCreateInfoNV = C.VkPipelineCoverageModulationStateCreateInfoNV

@[typedef]
pub struct C.VkPipelineCoverageModulationStateCreateInfoNV {
pub mut:
	sType                         StructureType = StructureType.pipeline_coverage_modulation_state_create_info_nv
	pNext                         voidptr       = unsafe { nil }
	flags                         PipelineCoverageModulationStateCreateFlagsNV
	coverageModulationMode        CoverageModulationModeNV
	coverageModulationTableEnable Bool32
	coverageModulationTableCount  u32
	pCoverageModulationTable      &f32
}

pub type AttachmentSampleCountInfoNV = C.VkAttachmentSampleCountInfoAMD

pub const nv_fill_rectangle_spec_version = 1
pub const nv_fill_rectangle_extension_name = c'VK_NV_fill_rectangle'

pub const nv_shader_sm_builtins_spec_version = 1
pub const nv_shader_sm_builtins_extension_name = c'VK_NV_shader_sm_builtins'
// PhysicalDeviceShaderSMBuiltinsPropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceShaderSMBuiltinsPropertiesNV = C.VkPhysicalDeviceShaderSMBuiltinsPropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceShaderSMBuiltinsPropertiesNV {
pub mut:
	sType            StructureType = StructureType.physical_device_shader_sm_builtins_properties_nv
	pNext            voidptr       = unsafe { nil }
	shaderSMCount    u32
	shaderWarpsPerSM u32
}

// PhysicalDeviceShaderSMBuiltinsFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderSMBuiltinsFeaturesNV = C.VkPhysicalDeviceShaderSMBuiltinsFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceShaderSMBuiltinsFeaturesNV {
pub mut:
	sType            StructureType = StructureType.physical_device_shader_sm_builtins_features_nv
	pNext            voidptr       = unsafe { nil }
	shaderSMBuiltins Bool32
}

pub const ext_post_depth_coverage_spec_version = 1
pub const ext_post_depth_coverage_extension_name = c'VK_EXT_post_depth_coverage'

pub const ext_image_drm_format_modifier_spec_version = 2
pub const ext_image_drm_format_modifier_extension_name = c'VK_EXT_image_drm_format_modifier'

pub type DrmFormatModifierPropertiesEXT = C.VkDrmFormatModifierPropertiesEXT

@[typedef]
pub struct C.VkDrmFormatModifierPropertiesEXT {
pub mut:
	drmFormatModifier               u64
	drmFormatModifierPlaneCount     u32
	drmFormatModifierTilingFeatures FormatFeatureFlags
}

// DrmFormatModifierPropertiesListEXT extends VkFormatProperties2
pub type DrmFormatModifierPropertiesListEXT = C.VkDrmFormatModifierPropertiesListEXT

@[typedef]
pub struct C.VkDrmFormatModifierPropertiesListEXT {
pub mut:
	sType                        StructureType = StructureType.drm_format_modifier_properties_list_ext
	pNext                        voidptr       = unsafe { nil }
	drmFormatModifierCount       u32
	pDrmFormatModifierProperties &DrmFormatModifierPropertiesEXT
}

// PhysicalDeviceImageDrmFormatModifierInfoEXT extends VkPhysicalDeviceImageFormatInfo2
pub type PhysicalDeviceImageDrmFormatModifierInfoEXT = C.VkPhysicalDeviceImageDrmFormatModifierInfoEXT

@[typedef]
pub struct C.VkPhysicalDeviceImageDrmFormatModifierInfoEXT {
pub mut:
	sType                 StructureType = StructureType.physical_device_image_drm_format_modifier_info_ext
	pNext                 voidptr       = unsafe { nil }
	drmFormatModifier     u64
	sharingMode           SharingMode
	queueFamilyIndexCount u32
	pQueueFamilyIndices   &u32
}

// ImageDrmFormatModifierListCreateInfoEXT extends VkImageCreateInfo
pub type ImageDrmFormatModifierListCreateInfoEXT = C.VkImageDrmFormatModifierListCreateInfoEXT

@[typedef]
pub struct C.VkImageDrmFormatModifierListCreateInfoEXT {
pub mut:
	sType                  StructureType = StructureType.image_drm_format_modifier_list_create_info_ext
	pNext                  voidptr       = unsafe { nil }
	drmFormatModifierCount u32
	pDrmFormatModifiers    &u64
}

// ImageDrmFormatModifierExplicitCreateInfoEXT extends VkImageCreateInfo
pub type ImageDrmFormatModifierExplicitCreateInfoEXT = C.VkImageDrmFormatModifierExplicitCreateInfoEXT

@[typedef]
pub struct C.VkImageDrmFormatModifierExplicitCreateInfoEXT {
pub mut:
	sType                       StructureType = StructureType.image_drm_format_modifier_explicit_create_info_ext
	pNext                       voidptr       = unsafe { nil }
	drmFormatModifier           u64
	drmFormatModifierPlaneCount u32
	pPlaneLayouts               &SubresourceLayout
}

pub type ImageDrmFormatModifierPropertiesEXT = C.VkImageDrmFormatModifierPropertiesEXT

@[typedef]
pub struct C.VkImageDrmFormatModifierPropertiesEXT {
pub mut:
	sType             StructureType = StructureType.image_drm_format_modifier_properties_ext
	pNext             voidptr       = unsafe { nil }
	drmFormatModifier u64
}

pub type DrmFormatModifierProperties2EXT = C.VkDrmFormatModifierProperties2EXT

@[typedef]
pub struct C.VkDrmFormatModifierProperties2EXT {
pub mut:
	drmFormatModifier               u64
	drmFormatModifierPlaneCount     u32
	drmFormatModifierTilingFeatures FormatFeatureFlags2
}

// DrmFormatModifierPropertiesList2EXT extends VkFormatProperties2
pub type DrmFormatModifierPropertiesList2EXT = C.VkDrmFormatModifierPropertiesList2EXT

@[typedef]
pub struct C.VkDrmFormatModifierPropertiesList2EXT {
pub mut:
	sType                        StructureType = StructureType.drm_format_modifier_properties_list2_ext
	pNext                        voidptr       = unsafe { nil }
	drmFormatModifierCount       u32
	pDrmFormatModifierProperties &DrmFormatModifierProperties2EXT
}

@[keep_args_alive]
fn C.vkGetImageDrmFormatModifierPropertiesEXT(device Device, image Image, mut p_properties ImageDrmFormatModifierPropertiesEXT) Result

pub type PFN_vkGetImageDrmFormatModifierPropertiesEXT = fn (device Device, image Image, mut p_properties ImageDrmFormatModifierPropertiesEXT) Result

@[inline]
pub fn get_image_drm_format_modifier_properties_ext(device Device,
	image Image,
	mut p_properties ImageDrmFormatModifierPropertiesEXT) Result {
	return C.vkGetImageDrmFormatModifierPropertiesEXT(device, image, mut p_properties)
}

// Pointer to VkValidationCacheEXT_T
pub type ValidationCacheEXT = voidptr

pub const ext_validation_cache_spec_version = 1
pub const ext_validation_cache_extension_name = c'VK_EXT_validation_cache'

pub enum ValidationCacheHeaderVersionEXT as u32 {
	one          = 1
	max_enum_ext = max_int
}
pub type ValidationCacheCreateFlagsEXT = u32
pub type ValidationCacheCreateInfoEXT = C.VkValidationCacheCreateInfoEXT

@[typedef]
pub struct C.VkValidationCacheCreateInfoEXT {
pub mut:
	sType           StructureType = StructureType.validation_cache_create_info_ext
	pNext           voidptr       = unsafe { nil }
	flags           ValidationCacheCreateFlagsEXT
	initialDataSize usize
	pInitialData    voidptr
}

// ShaderModuleValidationCacheCreateInfoEXT extends VkShaderModuleCreateInfo,VkPipelineShaderStageCreateInfo
pub type ShaderModuleValidationCacheCreateInfoEXT = C.VkShaderModuleValidationCacheCreateInfoEXT

@[typedef]
pub struct C.VkShaderModuleValidationCacheCreateInfoEXT {
pub mut:
	sType           StructureType = StructureType.shader_module_validation_cache_create_info_ext
	pNext           voidptr       = unsafe { nil }
	validationCache ValidationCacheEXT
}

@[keep_args_alive]
fn C.vkCreateValidationCacheEXT(device Device, p_create_info &ValidationCacheCreateInfoEXT, p_allocator &AllocationCallbacks, p_validation_cache &ValidationCacheEXT) Result

pub type PFN_vkCreateValidationCacheEXT = fn (device Device, p_create_info &ValidationCacheCreateInfoEXT, p_allocator &AllocationCallbacks, p_validation_cache &ValidationCacheEXT) Result

@[inline]
pub fn create_validation_cache_ext(device Device,
	p_create_info &ValidationCacheCreateInfoEXT,
	p_allocator &AllocationCallbacks,
	p_validation_cache &ValidationCacheEXT) Result {
	return C.vkCreateValidationCacheEXT(device, p_create_info, p_allocator, p_validation_cache)
}

@[keep_args_alive]
fn C.vkDestroyValidationCacheEXT(device Device, validation_cache ValidationCacheEXT, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyValidationCacheEXT = fn (device Device, validation_cache ValidationCacheEXT, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_validation_cache_ext(device Device,
	validation_cache ValidationCacheEXT,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyValidationCacheEXT(device, validation_cache, p_allocator)
}

@[keep_args_alive]
fn C.vkMergeValidationCachesEXT(device Device, dst_cache ValidationCacheEXT, src_cache_count u32, p_src_caches &ValidationCacheEXT) Result

pub type PFN_vkMergeValidationCachesEXT = fn (device Device, dst_cache ValidationCacheEXT, src_cache_count u32, p_src_caches &ValidationCacheEXT) Result

@[inline]
pub fn merge_validation_caches_ext(device Device,
	dst_cache ValidationCacheEXT,
	src_cache_count u32,
	p_src_caches &ValidationCacheEXT) Result {
	return C.vkMergeValidationCachesEXT(device, dst_cache, src_cache_count, p_src_caches)
}

@[keep_args_alive]
fn C.vkGetValidationCacheDataEXT(device Device, validation_cache ValidationCacheEXT, p_data_size &usize, p_data voidptr) Result

pub type PFN_vkGetValidationCacheDataEXT = fn (device Device, validation_cache ValidationCacheEXT, p_data_size &usize, p_data voidptr) Result

@[inline]
pub fn get_validation_cache_data_ext(device Device,
	validation_cache ValidationCacheEXT,
	p_data_size &usize,
	p_data voidptr) Result {
	return C.vkGetValidationCacheDataEXT(device, validation_cache, p_data_size, p_data)
}

pub const ext_descriptor_indexing_spec_version = 2
pub const ext_descriptor_indexing_extension_name = c'VK_EXT_descriptor_indexing'

pub type DescriptorBindingFlagBitsEXT = DescriptorBindingFlagBits

pub type DescriptorBindingFlagsEXT = u32
pub type DescriptorSetLayoutBindingFlagsCreateInfoEXT = C.VkDescriptorSetLayoutBindingFlagsCreateInfo

pub type PhysicalDeviceDescriptorIndexingFeaturesEXT = C.VkPhysicalDeviceDescriptorIndexingFeatures

pub type PhysicalDeviceDescriptorIndexingPropertiesEXT = C.VkPhysicalDeviceDescriptorIndexingProperties

pub type DescriptorSetVariableDescriptorCountAllocateInfoEXT = C.VkDescriptorSetVariableDescriptorCountAllocateInfo

pub type DescriptorSetVariableDescriptorCountLayoutSupportEXT = C.VkDescriptorSetVariableDescriptorCountLayoutSupport

pub const ext_shader_viewport_index_layer_spec_version = 1
pub const ext_shader_viewport_index_layer_extension_name = c'VK_EXT_shader_viewport_index_layer'

pub const nv_shading_rate_image_spec_version = 3
pub const nv_shading_rate_image_extension_name = c'VK_NV_shading_rate_image'

pub enum ShadingRatePaletteEntryNV as u32 {
	no_invocations              = 0
	_16_invocations_per_pixel   = 1
	_8_invocations_per_pixel    = 2
	_4_invocations_per_pixel    = 3
	_2_invocations_per_pixel    = 4
	_1_invocation_per_pixel     = 5
	_1_invocation_per2x1_pixels = 6
	_1_invocation_per1x2_pixels = 7
	_1_invocation_per2x2_pixels = 8
	_1_invocation_per4x2_pixels = 9
	_1_invocation_per2x4_pixels = 10
	_1_invocation_per4x4_pixels = 11
	max_enum_nv                 = max_int
}

pub enum CoarseSampleOrderTypeNV as u32 {
	default      = 0
	custom       = 1
	pixel_major  = 2
	sample_major = 3
	max_enum_nv  = max_int
}
pub type ShadingRatePaletteNV = C.VkShadingRatePaletteNV

@[typedef]
pub struct C.VkShadingRatePaletteNV {
pub mut:
	shadingRatePaletteEntryCount u32
	pShadingRatePaletteEntries   &ShadingRatePaletteEntryNV
}

// PipelineViewportShadingRateImageStateCreateInfoNV extends VkPipelineViewportStateCreateInfo
pub type PipelineViewportShadingRateImageStateCreateInfoNV = C.VkPipelineViewportShadingRateImageStateCreateInfoNV

@[typedef]
pub struct C.VkPipelineViewportShadingRateImageStateCreateInfoNV {
pub mut:
	sType                  StructureType = StructureType.pipeline_viewport_shading_rate_image_state_create_info_nv
	pNext                  voidptr       = unsafe { nil }
	shadingRateImageEnable Bool32
	viewportCount          u32
	pShadingRatePalettes   &ShadingRatePaletteNV
}

// PhysicalDeviceShadingRateImageFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShadingRateImageFeaturesNV = C.VkPhysicalDeviceShadingRateImageFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceShadingRateImageFeaturesNV {
pub mut:
	sType                        StructureType = StructureType.physical_device_shading_rate_image_features_nv
	pNext                        voidptr       = unsafe { nil }
	shadingRateImage             Bool32
	shadingRateCoarseSampleOrder Bool32
}

// PhysicalDeviceShadingRateImagePropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceShadingRateImagePropertiesNV = C.VkPhysicalDeviceShadingRateImagePropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceShadingRateImagePropertiesNV {
pub mut:
	sType                       StructureType = StructureType.physical_device_shading_rate_image_properties_nv
	pNext                       voidptr       = unsafe { nil }
	shadingRateTexelSize        Extent2D
	shadingRatePaletteSize      u32
	shadingRateMaxCoarseSamples u32
}

pub type CoarseSampleLocationNV = C.VkCoarseSampleLocationNV

@[typedef]
pub struct C.VkCoarseSampleLocationNV {
pub mut:
	pixelX u32
	pixelY u32
	sample u32
}

pub type CoarseSampleOrderCustomNV = C.VkCoarseSampleOrderCustomNV

@[typedef]
pub struct C.VkCoarseSampleOrderCustomNV {
pub mut:
	shadingRate         ShadingRatePaletteEntryNV
	sampleCount         u32
	sampleLocationCount u32
	pSampleLocations    &CoarseSampleLocationNV
}

// PipelineViewportCoarseSampleOrderStateCreateInfoNV extends VkPipelineViewportStateCreateInfo
pub type PipelineViewportCoarseSampleOrderStateCreateInfoNV = C.VkPipelineViewportCoarseSampleOrderStateCreateInfoNV

@[typedef]
pub struct C.VkPipelineViewportCoarseSampleOrderStateCreateInfoNV {
pub mut:
	sType                  StructureType = StructureType.pipeline_viewport_coarse_sample_order_state_create_info_nv
	pNext                  voidptr       = unsafe { nil }
	sampleOrderType        CoarseSampleOrderTypeNV
	customSampleOrderCount u32
	pCustomSampleOrders    &CoarseSampleOrderCustomNV
}

@[keep_args_alive]
fn C.vkCmdBindShadingRateImageNV(command_buffer CommandBuffer, image_view ImageView, image_layout ImageLayout)

pub type PFN_vkCmdBindShadingRateImageNV = fn (command_buffer CommandBuffer, image_view ImageView, image_layout ImageLayout)

@[inline]
pub fn cmd_bind_shading_rate_image_nv(command_buffer CommandBuffer,
	image_view ImageView,
	image_layout ImageLayout) {
	C.vkCmdBindShadingRateImageNV(command_buffer, image_view, image_layout)
}

@[keep_args_alive]
fn C.vkCmdSetViewportShadingRatePaletteNV(command_buffer CommandBuffer, first_viewport u32, viewport_count u32, p_shading_rate_palettes &ShadingRatePaletteNV)

pub type PFN_vkCmdSetViewportShadingRatePaletteNV = fn (command_buffer CommandBuffer, first_viewport u32, viewport_count u32, p_shading_rate_palettes &ShadingRatePaletteNV)

@[inline]
pub fn cmd_set_viewport_shading_rate_palette_nv(command_buffer CommandBuffer,
	first_viewport u32,
	viewport_count u32,
	p_shading_rate_palettes &ShadingRatePaletteNV) {
	C.vkCmdSetViewportShadingRatePaletteNV(command_buffer, first_viewport, viewport_count,
		p_shading_rate_palettes)
}

@[keep_args_alive]
fn C.vkCmdSetCoarseSampleOrderNV(command_buffer CommandBuffer, sample_order_type CoarseSampleOrderTypeNV, custom_sample_order_count u32, p_custom_sample_orders &CoarseSampleOrderCustomNV)

pub type PFN_vkCmdSetCoarseSampleOrderNV = fn (command_buffer CommandBuffer, sample_order_type CoarseSampleOrderTypeNV, custom_sample_order_count u32, p_custom_sample_orders &CoarseSampleOrderCustomNV)

@[inline]
pub fn cmd_set_coarse_sample_order_nv(command_buffer CommandBuffer,
	sample_order_type CoarseSampleOrderTypeNV,
	custom_sample_order_count u32,
	p_custom_sample_orders &CoarseSampleOrderCustomNV) {
	C.vkCmdSetCoarseSampleOrderNV(command_buffer, sample_order_type, custom_sample_order_count,
		p_custom_sample_orders)
}

// Pointer to VkAccelerationStructureNV_T
pub type AccelerationStructureNV = voidptr

pub const nv_ray_tracing_spec_version = 3
pub const nv_ray_tracing_extension_name = c'VK_NV_ray_tracing'
pub const shader_unused_khr = ~u32(0)
pub const shader_unused_nv = shader_unused_khr

pub enum RayTracingShaderGroupTypeKHR as u32 {
	general              = 0
	triangles_hit_group  = 1
	procedural_hit_group = 2
	max_enum_khr         = max_int
}
pub type RayTracingShaderGroupTypeNV = RayTracingShaderGroupTypeKHR

pub enum GeometryTypeKHR as u32 {
	triangles               = 0
	aabbs                   = 1
	instances               = 2
	spheres_nv              = 1000429004
	linear_swept_spheres_nv = 1000429005
	max_enum_khr            = max_int
}
pub type GeometryTypeNV = GeometryTypeKHR

pub enum AccelerationStructureTypeKHR as u32 {
	top_level    = 0
	bottom_level = 1
	generic      = 2
	max_enum_khr = max_int
}
pub type AccelerationStructureTypeNV = AccelerationStructureTypeKHR

pub enum CopyAccelerationStructureModeKHR as u32 {
	clone        = 0
	compact      = 1
	serialize    = 2
	deserialize  = 3
	max_enum_khr = max_int
}
pub type CopyAccelerationStructureModeNV = CopyAccelerationStructureModeKHR

pub enum AccelerationStructureMemoryRequirementsTypeNV as u32 {
	object         = 0
	build_scratch  = 1
	update_scratch = 2
	max_enum_nv    = max_int
}

pub enum GeometryFlagBitsKHR as u32 {
	opaque                          = u32(0x00000001)
	no_duplicate_any_hit_invocation = u32(0x00000002)
	max_enum_khr                    = max_int
}
pub type GeometryFlagsKHR = u32
pub type GeometryFlagsNV = u32
pub type GeometryFlagBitsNV = GeometryFlagBitsKHR

pub enum GeometryInstanceFlagBitsKHR as u32 {
	triangle_facing_cull_disable          = u32(0x00000001)
	triangle_flip_facing                  = u32(0x00000002)
	force_opaque                          = u32(0x00000004)
	force_no_opaque                       = u32(0x00000008)
	force_opacity_micromap2_state_bit_ext = u32(0x00000010)
	disable_opacity_micromaps_bit_ext     = u32(0x00000020)
	max_enum_khr                          = max_int
}
pub type GeometryInstanceFlagsKHR = u32
pub type GeometryInstanceFlagsNV = u32
pub type GeometryInstanceFlagBitsNV = GeometryInstanceFlagBitsKHR

pub enum BuildAccelerationStructureFlagBitsKHR as u32 {
	allow_update                               = u32(0x00000001)
	allow_compaction                           = u32(0x00000002)
	prefer_fast_trace                          = u32(0x00000004)
	prefer_fast_build                          = u32(0x00000008)
	low_memory                                 = u32(0x00000010)
	motion_bit_nv                              = u32(0x00000020)
	allow_opacity_micromap_update_bit_ext      = u32(0x00000040)
	allow_disable_opacity_micromaps_bit_ext    = u32(0x00000080)
	allow_opacity_micromap_data_update_bit_ext = u32(0x00000100)
	allow_data_access                          = u32(0x00000800)
	allow_cluster_opacity_micromaps_bit_nv     = u32(0x00001000)
	max_enum_khr                               = max_int
}
pub type BuildAccelerationStructureFlagsKHR = u32
pub type BuildAccelerationStructureFlagsNV = u32
pub type BuildAccelerationStructureFlagBitsNV = BuildAccelerationStructureFlagBitsKHR

pub type RayTracingShaderGroupCreateInfoNV = C.VkRayTracingShaderGroupCreateInfoNV

@[typedef]
pub struct C.VkRayTracingShaderGroupCreateInfoNV {
pub mut:
	sType              StructureType = StructureType.ray_tracing_shader_group_create_info_nv
	pNext              voidptr       = unsafe { nil }
	type               RayTracingShaderGroupTypeKHR
	generalShader      u32
	closestHitShader   u32
	anyHitShader       u32
	intersectionShader u32
}

pub type RayTracingPipelineCreateInfoNV = C.VkRayTracingPipelineCreateInfoNV

@[typedef]
pub struct C.VkRayTracingPipelineCreateInfoNV {
pub mut:
	sType              StructureType = StructureType.ray_tracing_pipeline_create_info_nv
	pNext              voidptr       = unsafe { nil }
	flags              PipelineCreateFlags
	stageCount         u32
	pStages            &PipelineShaderStageCreateInfo
	groupCount         u32
	pGroups            &RayTracingShaderGroupCreateInfoNV
	maxRecursionDepth  u32
	layout             PipelineLayout
	basePipelineHandle Pipeline
	basePipelineIndex  i32
}

pub type GeometryTrianglesNV = C.VkGeometryTrianglesNV

@[typedef]
pub struct C.VkGeometryTrianglesNV {
pub mut:
	sType           StructureType = StructureType.geometry_triangles_nv
	pNext           voidptr       = unsafe { nil }
	vertexData      Buffer
	vertexOffset    DeviceSize
	vertexCount     u32
	vertexStride    DeviceSize
	vertexFormat    Format
	indexData       Buffer
	indexOffset     DeviceSize
	indexCount      u32
	indexType       IndexType
	transformData   Buffer
	transformOffset DeviceSize
}

pub type GeometryAABBNV = C.VkGeometryAABBNV

@[typedef]
pub struct C.VkGeometryAABBNV {
pub mut:
	sType    StructureType = StructureType.geometry_aabb_nv
	pNext    voidptr       = unsafe { nil }
	aabbData Buffer
	numAABBs u32
	stride   u32
	offset   DeviceSize
}

pub type GeometryDataNV = C.VkGeometryDataNV

@[typedef]
pub struct C.VkGeometryDataNV {
pub mut:
	triangles GeometryTrianglesNV
	aabbs     GeometryAABBNV
}

pub type GeometryNV = C.VkGeometryNV

@[typedef]
pub struct C.VkGeometryNV {
pub mut:
	sType        StructureType = StructureType.geometry_nv
	pNext        voidptr       = unsafe { nil }
	geometryType GeometryTypeKHR
	geometry     GeometryDataNV
	flags        GeometryFlagsKHR
}

pub type AccelerationStructureInfoNV = C.VkAccelerationStructureInfoNV

@[typedef]
pub struct C.VkAccelerationStructureInfoNV {
pub mut:
	sType         StructureType = StructureType.acceleration_structure_info_nv
	pNext         voidptr       = unsafe { nil }
	type          AccelerationStructureTypeNV
	flags         BuildAccelerationStructureFlagsNV
	instanceCount u32
	geometryCount u32
	pGeometries   &GeometryNV
}

pub type AccelerationStructureCreateInfoNV = C.VkAccelerationStructureCreateInfoNV

@[typedef]
pub struct C.VkAccelerationStructureCreateInfoNV {
pub mut:
	sType         StructureType = StructureType.acceleration_structure_create_info_nv
	pNext         voidptr       = unsafe { nil }
	compactedSize DeviceSize
	info          AccelerationStructureInfoNV
}

pub type BindAccelerationStructureMemoryInfoNV = C.VkBindAccelerationStructureMemoryInfoNV

@[typedef]
pub struct C.VkBindAccelerationStructureMemoryInfoNV {
pub mut:
	sType                 StructureType = StructureType.bind_acceleration_structure_memory_info_nv
	pNext                 voidptr       = unsafe { nil }
	accelerationStructure AccelerationStructureNV
	memory                DeviceMemory
	memoryOffset          DeviceSize
	deviceIndexCount      u32
	pDeviceIndices        &u32
}

// WriteDescriptorSetAccelerationStructureNV extends VkWriteDescriptorSet
pub type WriteDescriptorSetAccelerationStructureNV = C.VkWriteDescriptorSetAccelerationStructureNV

@[typedef]
pub struct C.VkWriteDescriptorSetAccelerationStructureNV {
pub mut:
	sType                      StructureType = StructureType.write_descriptor_set_acceleration_structure_nv
	pNext                      voidptr       = unsafe { nil }
	accelerationStructureCount u32
	pAccelerationStructures    &AccelerationStructureNV
}

pub type AccelerationStructureMemoryRequirementsInfoNV = C.VkAccelerationStructureMemoryRequirementsInfoNV

@[typedef]
pub struct C.VkAccelerationStructureMemoryRequirementsInfoNV {
pub mut:
	sType                 StructureType = StructureType.acceleration_structure_memory_requirements_info_nv
	pNext                 voidptr       = unsafe { nil }
	type                  AccelerationStructureMemoryRequirementsTypeNV
	accelerationStructure AccelerationStructureNV
}

// PhysicalDeviceRayTracingPropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceRayTracingPropertiesNV = C.VkPhysicalDeviceRayTracingPropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceRayTracingPropertiesNV {
pub mut:
	sType                                  StructureType = StructureType.physical_device_ray_tracing_properties_nv
	pNext                                  voidptr       = unsafe { nil }
	shaderGroupHandleSize                  u32
	maxRecursionDepth                      u32
	maxShaderGroupStride                   u32
	shaderGroupBaseAlignment               u32
	maxGeometryCount                       u64
	maxInstanceCount                       u64
	maxTriangleCount                       u64
	maxDescriptorSetAccelerationStructures u32
}

pub type TransformMatrixKHR = C.VkTransformMatrixKHR

@[typedef]
pub struct C.VkTransformMatrixKHR {
pub mut:
	matrix [4][3]f32
}

pub type TransformMatrixNV = C.VkTransformMatrixKHR

pub type AabbPositionsKHR = C.VkAabbPositionsKHR

@[typedef]
pub struct C.VkAabbPositionsKHR {
pub mut:
	minX f32
	minY f32
	minZ f32
	maxX f32
	maxY f32
	maxZ f32
}

pub type AabbPositionsNV = C.VkAabbPositionsKHR

pub type AccelerationStructureInstanceKHR = C.VkAccelerationStructureInstanceKHR

@[typedef]
pub struct C.VkAccelerationStructureInstanceKHR {
pub mut:
	transform                              TransformMatrixKHR
	instanceCustomIndex                    u32
	mask                                   u32
	instanceShaderBindingTableRecordOffset u32
	flags                                  GeometryInstanceFlagsKHR
	accelerationStructureReference         u64
}

pub type AccelerationStructureInstanceNV = C.VkAccelerationStructureInstanceKHR

@[keep_args_alive]
fn C.vkCreateAccelerationStructureNV(device Device, p_create_info &AccelerationStructureCreateInfoNV, p_allocator &AllocationCallbacks, p_acceleration_structure &AccelerationStructureNV) Result

pub type PFN_vkCreateAccelerationStructureNV = fn (device Device, p_create_info &AccelerationStructureCreateInfoNV, p_allocator &AllocationCallbacks, p_acceleration_structure &AccelerationStructureNV) Result

@[inline]
pub fn create_acceleration_structure_nv(device Device,
	p_create_info &AccelerationStructureCreateInfoNV,
	p_allocator &AllocationCallbacks,
	p_acceleration_structure &AccelerationStructureNV) Result {
	return C.vkCreateAccelerationStructureNV(device, p_create_info, p_allocator, p_acceleration_structure)
}

@[keep_args_alive]
fn C.vkDestroyAccelerationStructureNV(device Device, acceleration_structure AccelerationStructureNV, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyAccelerationStructureNV = fn (device Device, acceleration_structure AccelerationStructureNV, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_acceleration_structure_nv(device Device,
	acceleration_structure AccelerationStructureNV,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyAccelerationStructureNV(device, acceleration_structure, p_allocator)
}

@[keep_args_alive]
fn C.vkGetAccelerationStructureMemoryRequirementsNV(device Device, p_info &AccelerationStructureMemoryRequirementsInfoNV, mut p_memory_requirements MemoryRequirements2KHR)

pub type PFN_vkGetAccelerationStructureMemoryRequirementsNV = fn (device Device, p_info &AccelerationStructureMemoryRequirementsInfoNV, mut p_memory_requirements MemoryRequirements2KHR)

@[inline]
pub fn get_acceleration_structure_memory_requirements_nv(device Device,
	p_info &AccelerationStructureMemoryRequirementsInfoNV,
	mut p_memory_requirements MemoryRequirements2KHR) {
	C.vkGetAccelerationStructureMemoryRequirementsNV(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkBindAccelerationStructureMemoryNV(device Device, bind_info_count u32, p_bind_infos &BindAccelerationStructureMemoryInfoNV) Result

pub type PFN_vkBindAccelerationStructureMemoryNV = fn (device Device, bind_info_count u32, p_bind_infos &BindAccelerationStructureMemoryInfoNV) Result

@[inline]
pub fn bind_acceleration_structure_memory_nv(device Device,
	bind_info_count u32,
	p_bind_infos &BindAccelerationStructureMemoryInfoNV) Result {
	return C.vkBindAccelerationStructureMemoryNV(device, bind_info_count, p_bind_infos)
}

@[keep_args_alive]
fn C.vkCmdBuildAccelerationStructureNV(command_buffer CommandBuffer, p_info &AccelerationStructureInfoNV, instance_data Buffer, instance_offset DeviceSize, update Bool32, dst AccelerationStructureNV, src AccelerationStructureNV, scratch Buffer, scratch_offset DeviceSize)

pub type PFN_vkCmdBuildAccelerationStructureNV = fn (command_buffer CommandBuffer, p_info &AccelerationStructureInfoNV, instance_data Buffer, instance_offset DeviceSize, update Bool32, dst AccelerationStructureNV, src AccelerationStructureNV, scratch Buffer, scratch_offset DeviceSize)

@[inline]
pub fn cmd_build_acceleration_structure_nv(command_buffer CommandBuffer,
	p_info &AccelerationStructureInfoNV,
	instance_data Buffer,
	instance_offset DeviceSize,
	update Bool32,
	dst AccelerationStructureNV,
	src AccelerationStructureNV,
	scratch Buffer,
	scratch_offset DeviceSize) {
	C.vkCmdBuildAccelerationStructureNV(command_buffer, p_info, instance_data, instance_offset,
		update, dst, src, scratch, scratch_offset)
}

@[keep_args_alive]
fn C.vkCmdCopyAccelerationStructureNV(command_buffer CommandBuffer, dst AccelerationStructureNV, src AccelerationStructureNV, mode CopyAccelerationStructureModeKHR)

pub type PFN_vkCmdCopyAccelerationStructureNV = fn (command_buffer CommandBuffer, dst AccelerationStructureNV, src AccelerationStructureNV, mode CopyAccelerationStructureModeKHR)

@[inline]
pub fn cmd_copy_acceleration_structure_nv(command_buffer CommandBuffer,
	dst AccelerationStructureNV,
	src AccelerationStructureNV,
	mode CopyAccelerationStructureModeKHR) {
	C.vkCmdCopyAccelerationStructureNV(command_buffer, dst, src, mode)
}

@[keep_args_alive]
fn C.vkCmdTraceRaysNV(command_buffer CommandBuffer, raygen_shader_binding_table_buffer Buffer, raygen_shader_binding_offset DeviceSize, miss_shader_binding_table_buffer Buffer, miss_shader_binding_offset DeviceSize, miss_shader_binding_stride DeviceSize, hit_shader_binding_table_buffer Buffer, hit_shader_binding_offset DeviceSize, hit_shader_binding_stride DeviceSize, callable_shader_binding_table_buffer Buffer, callable_shader_binding_offset DeviceSize, callable_shader_binding_stride DeviceSize, width u32, height u32, depth u32)

pub type PFN_vkCmdTraceRaysNV = fn (command_buffer CommandBuffer, raygen_shader_binding_table_buffer Buffer, raygen_shader_binding_offset DeviceSize, miss_shader_binding_table_buffer Buffer, miss_shader_binding_offset DeviceSize, miss_shader_binding_stride DeviceSize, hit_shader_binding_table_buffer Buffer, hit_shader_binding_offset DeviceSize, hit_shader_binding_stride DeviceSize, callable_shader_binding_table_buffer Buffer, callable_shader_binding_offset DeviceSize, callable_shader_binding_stride DeviceSize, width u32, height u32, depth u32)

@[inline]
pub fn cmd_trace_rays_nv(command_buffer CommandBuffer,
	raygen_shader_binding_table_buffer Buffer,
	raygen_shader_binding_offset DeviceSize,
	miss_shader_binding_table_buffer Buffer,
	miss_shader_binding_offset DeviceSize,
	miss_shader_binding_stride DeviceSize,
	hit_shader_binding_table_buffer Buffer,
	hit_shader_binding_offset DeviceSize,
	hit_shader_binding_stride DeviceSize,
	callable_shader_binding_table_buffer Buffer,
	callable_shader_binding_offset DeviceSize,
	callable_shader_binding_stride DeviceSize,
	width u32,
	height u32,
	depth u32) {
	C.vkCmdTraceRaysNV(command_buffer, raygen_shader_binding_table_buffer, raygen_shader_binding_offset,
		miss_shader_binding_table_buffer, miss_shader_binding_offset, miss_shader_binding_stride,
		hit_shader_binding_table_buffer, hit_shader_binding_offset, hit_shader_binding_stride,
		callable_shader_binding_table_buffer, callable_shader_binding_offset, callable_shader_binding_stride,
		width, height, depth)
}

@[keep_args_alive]
fn C.vkCreateRayTracingPipelinesNV(device Device, pipeline_cache PipelineCache, create_info_count u32, p_create_infos &RayTracingPipelineCreateInfoNV, p_allocator &AllocationCallbacks, p_pipelines &Pipeline) Result

pub type PFN_vkCreateRayTracingPipelinesNV = fn (device Device, pipeline_cache PipelineCache, create_info_count u32, p_create_infos &RayTracingPipelineCreateInfoNV, p_allocator &AllocationCallbacks, p_pipelines &Pipeline) Result

@[inline]
pub fn create_ray_tracing_pipelines_nv(device Device,
	pipeline_cache PipelineCache,
	create_info_count u32,
	p_create_infos &RayTracingPipelineCreateInfoNV,
	p_allocator &AllocationCallbacks,
	p_pipelines &Pipeline) Result {
	return C.vkCreateRayTracingPipelinesNV(device, pipeline_cache, create_info_count,
		p_create_infos, p_allocator, p_pipelines)
}

@[keep_args_alive]
fn C.vkGetRayTracingShaderGroupHandlesKHR(device Device, pipeline Pipeline, first_group u32, group_count u32, data_size usize, p_data voidptr) Result

pub type PFN_vkGetRayTracingShaderGroupHandlesKHR = fn (device Device, pipeline Pipeline, first_group u32, group_count u32, data_size usize, p_data voidptr) Result

@[inline]
pub fn get_ray_tracing_shader_group_handles_khr(device Device,
	pipeline Pipeline,
	first_group u32,
	group_count u32,
	data_size usize,
	p_data voidptr) Result {
	return C.vkGetRayTracingShaderGroupHandlesKHR(device, pipeline, first_group, group_count,
		data_size, p_data)
}

@[keep_args_alive]
fn C.vkGetRayTracingShaderGroupHandlesNV(device Device, pipeline Pipeline, first_group u32, group_count u32, data_size usize, p_data voidptr) Result

pub type PFN_vkGetRayTracingShaderGroupHandlesNV = fn (device Device, pipeline Pipeline, first_group u32, group_count u32, data_size usize, p_data voidptr) Result

@[inline]
pub fn get_ray_tracing_shader_group_handles_nv(device Device,
	pipeline Pipeline,
	first_group u32,
	group_count u32,
	data_size usize,
	p_data voidptr) Result {
	return C.vkGetRayTracingShaderGroupHandlesNV(device, pipeline, first_group, group_count,
		data_size, p_data)
}

@[keep_args_alive]
fn C.vkGetAccelerationStructureHandleNV(device Device, acceleration_structure AccelerationStructureNV, data_size usize, p_data voidptr) Result

pub type PFN_vkGetAccelerationStructureHandleNV = fn (device Device, acceleration_structure AccelerationStructureNV, data_size usize, p_data voidptr) Result

@[inline]
pub fn get_acceleration_structure_handle_nv(device Device,
	acceleration_structure AccelerationStructureNV,
	data_size usize,
	p_data voidptr) Result {
	return C.vkGetAccelerationStructureHandleNV(device, acceleration_structure, data_size,
		p_data)
}

@[keep_args_alive]
fn C.vkCmdWriteAccelerationStructuresPropertiesNV(command_buffer CommandBuffer, acceleration_structure_count u32, p_acceleration_structures &AccelerationStructureNV, query_type QueryType, query_pool QueryPool, first_query u32)

pub type PFN_vkCmdWriteAccelerationStructuresPropertiesNV = fn (command_buffer CommandBuffer, acceleration_structure_count u32, p_acceleration_structures &AccelerationStructureNV, query_type QueryType, query_pool QueryPool, first_query u32)

@[inline]
pub fn cmd_write_acceleration_structures_properties_nv(command_buffer CommandBuffer,
	acceleration_structure_count u32,
	p_acceleration_structures &AccelerationStructureNV,
	query_type QueryType,
	query_pool QueryPool,
	first_query u32) {
	C.vkCmdWriteAccelerationStructuresPropertiesNV(command_buffer, acceleration_structure_count,
		p_acceleration_structures, query_type, query_pool, first_query)
}

@[keep_args_alive]
fn C.vkCompileDeferredNV(device Device, pipeline Pipeline, shader u32) Result

pub type PFN_vkCompileDeferredNV = fn (device Device, pipeline Pipeline, shader u32) Result

@[inline]
pub fn compile_deferred_nv(device Device,
	pipeline Pipeline,
	shader u32) Result {
	return C.vkCompileDeferredNV(device, pipeline, shader)
}

pub const nv_representative_fragment_test_spec_version = 2
pub const nv_representative_fragment_test_extension_name = c'VK_NV_representative_fragment_test'
// PhysicalDeviceRepresentativeFragmentTestFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRepresentativeFragmentTestFeaturesNV = C.VkPhysicalDeviceRepresentativeFragmentTestFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceRepresentativeFragmentTestFeaturesNV {
pub mut:
	sType                      StructureType = StructureType.physical_device_representative_fragment_test_features_nv
	pNext                      voidptr       = unsafe { nil }
	representativeFragmentTest Bool32
}

// PipelineRepresentativeFragmentTestStateCreateInfoNV extends VkGraphicsPipelineCreateInfo
pub type PipelineRepresentativeFragmentTestStateCreateInfoNV = C.VkPipelineRepresentativeFragmentTestStateCreateInfoNV

@[typedef]
pub struct C.VkPipelineRepresentativeFragmentTestStateCreateInfoNV {
pub mut:
	sType                            StructureType = StructureType.pipeline_representative_fragment_test_state_create_info_nv
	pNext                            voidptr       = unsafe { nil }
	representativeFragmentTestEnable Bool32
}

pub const ext_filter_cubic_spec_version = 3
pub const ext_filter_cubic_extension_name = c'VK_EXT_filter_cubic'
// PhysicalDeviceImageViewImageFormatInfoEXT extends VkPhysicalDeviceImageFormatInfo2
pub type PhysicalDeviceImageViewImageFormatInfoEXT = C.VkPhysicalDeviceImageViewImageFormatInfoEXT

@[typedef]
pub struct C.VkPhysicalDeviceImageViewImageFormatInfoEXT {
pub mut:
	sType         StructureType = StructureType.physical_device_image_view_image_format_info_ext
	pNext         voidptr       = unsafe { nil }
	imageViewType ImageViewType
}

// FilterCubicImageViewImageFormatPropertiesEXT extends VkImageFormatProperties2
pub type FilterCubicImageViewImageFormatPropertiesEXT = C.VkFilterCubicImageViewImageFormatPropertiesEXT

@[typedef]
pub struct C.VkFilterCubicImageViewImageFormatPropertiesEXT {
pub mut:
	sType             StructureType = StructureType.filter_cubic_image_view_image_format_properties_ext
	pNext             voidptr       = unsafe { nil }
	filterCubic       Bool32
	filterCubicMinmax Bool32
}

pub const qcom_render_pass_shader_resolve_spec_version = 4
pub const qcom_render_pass_shader_resolve_extension_name = c'VK_QCOM_render_pass_shader_resolve'

pub const ext_global_priority_spec_version = 2
pub const ext_global_priority_extension_name = c'VK_EXT_global_priority'

pub type QueueGlobalPriorityEXT = QueueGlobalPriority

pub type DeviceQueueGlobalPriorityCreateInfoEXT = C.VkDeviceQueueGlobalPriorityCreateInfo

pub const ext_external_memory_host_spec_version = 1
pub const ext_external_memory_host_extension_name = c'VK_EXT_external_memory_host'
// ImportMemoryHostPointerInfoEXT extends VkMemoryAllocateInfo
pub type ImportMemoryHostPointerInfoEXT = C.VkImportMemoryHostPointerInfoEXT

@[typedef]
pub struct C.VkImportMemoryHostPointerInfoEXT {
pub mut:
	sType        StructureType = StructureType.import_memory_host_pointer_info_ext
	pNext        voidptr       = unsafe { nil }
	handleType   ExternalMemoryHandleTypeFlagBits
	pHostPointer voidptr
}

pub type MemoryHostPointerPropertiesEXT = C.VkMemoryHostPointerPropertiesEXT

@[typedef]
pub struct C.VkMemoryHostPointerPropertiesEXT {
pub mut:
	sType          StructureType = StructureType.memory_host_pointer_properties_ext
	pNext          voidptr       = unsafe { nil }
	memoryTypeBits u32
}

// PhysicalDeviceExternalMemoryHostPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceExternalMemoryHostPropertiesEXT = C.VkPhysicalDeviceExternalMemoryHostPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceExternalMemoryHostPropertiesEXT {
pub mut:
	sType                           StructureType = StructureType.physical_device_external_memory_host_properties_ext
	pNext                           voidptr       = unsafe { nil }
	minImportedHostPointerAlignment DeviceSize
}

@[keep_args_alive]
fn C.vkGetMemoryHostPointerPropertiesEXT(device Device, handle_type ExternalMemoryHandleTypeFlagBits, p_host_pointer voidptr, mut p_memory_host_pointer_properties MemoryHostPointerPropertiesEXT) Result

pub type PFN_vkGetMemoryHostPointerPropertiesEXT = fn (device Device, handle_type ExternalMemoryHandleTypeFlagBits, p_host_pointer voidptr, mut p_memory_host_pointer_properties MemoryHostPointerPropertiesEXT) Result

@[inline]
pub fn get_memory_host_pointer_properties_ext(device Device,
	handle_type ExternalMemoryHandleTypeFlagBits,
	p_host_pointer voidptr,
	mut p_memory_host_pointer_properties MemoryHostPointerPropertiesEXT) Result {
	return C.vkGetMemoryHostPointerPropertiesEXT(device, handle_type, p_host_pointer, mut
		p_memory_host_pointer_properties)
}

pub const amd_buffer_marker_spec_version = 1
pub const amd_buffer_marker_extension_name = c'VK_AMD_buffer_marker'

@[keep_args_alive]
fn C.vkCmdWriteBufferMarkerAMD(command_buffer CommandBuffer, pipeline_stage PipelineStageFlagBits, dst_buffer Buffer, dst_offset DeviceSize, marker u32)

pub type PFN_vkCmdWriteBufferMarkerAMD = fn (command_buffer CommandBuffer, pipeline_stage PipelineStageFlagBits, dst_buffer Buffer, dst_offset DeviceSize, marker u32)

@[inline]
pub fn cmd_write_buffer_marker_amd(command_buffer CommandBuffer,
	pipeline_stage PipelineStageFlagBits,
	dst_buffer Buffer,
	dst_offset DeviceSize,
	marker u32) {
	C.vkCmdWriteBufferMarkerAMD(command_buffer, pipeline_stage, dst_buffer, dst_offset,
		marker)
}

@[keep_args_alive]
fn C.vkCmdWriteBufferMarker2AMD(command_buffer CommandBuffer, stage PipelineStageFlags2, dst_buffer Buffer, dst_offset DeviceSize, marker u32)

pub type PFN_vkCmdWriteBufferMarker2AMD = fn (command_buffer CommandBuffer, stage PipelineStageFlags2, dst_buffer Buffer, dst_offset DeviceSize, marker u32)

@[inline]
pub fn cmd_write_buffer_marker2_amd(command_buffer CommandBuffer,
	stage PipelineStageFlags2,
	dst_buffer Buffer,
	dst_offset DeviceSize,
	marker u32) {
	C.vkCmdWriteBufferMarker2AMD(command_buffer, stage, dst_buffer, dst_offset, marker)
}

pub const amd_pipeline_compiler_control_spec_version = 1
pub const amd_pipeline_compiler_control_extension_name = c'VK_AMD_pipeline_compiler_control'

pub enum PipelineCompilerControlFlagBitsAMD as u32 {
	max_enum_amd = max_int
}
pub type PipelineCompilerControlFlagsAMD = u32

// PipelineCompilerControlCreateInfoAMD extends VkGraphicsPipelineCreateInfo,VkComputePipelineCreateInfo
pub type PipelineCompilerControlCreateInfoAMD = C.VkPipelineCompilerControlCreateInfoAMD

@[typedef]
pub struct C.VkPipelineCompilerControlCreateInfoAMD {
pub mut:
	sType                StructureType = StructureType.pipeline_compiler_control_create_info_amd
	pNext                voidptr       = unsafe { nil }
	compilerControlFlags PipelineCompilerControlFlagsAMD
}

pub const ext_calibrated_timestamps_spec_version = 2
pub const ext_calibrated_timestamps_extension_name = c'VK_EXT_calibrated_timestamps'

pub type TimeDomainEXT = TimeDomainKHR

pub type CalibratedTimestampInfoEXT = C.VkCalibratedTimestampInfoKHR

@[keep_args_alive]
fn C.vkGetPhysicalDeviceCalibrateableTimeDomainsEXT(physical_device PhysicalDevice, p_time_domain_count &u32, p_time_domains &TimeDomainKHR) Result

pub type PFN_vkGetPhysicalDeviceCalibrateableTimeDomainsEXT = fn (physical_device PhysicalDevice, p_time_domain_count &u32, p_time_domains &TimeDomainKHR) Result

@[inline]
pub fn get_physical_device_calibrateable_time_domains_ext(physical_device PhysicalDevice,
	p_time_domain_count &u32,
	p_time_domains &TimeDomainKHR) Result {
	return C.vkGetPhysicalDeviceCalibrateableTimeDomainsEXT(physical_device, p_time_domain_count,
		p_time_domains)
}

@[keep_args_alive]
fn C.vkGetCalibratedTimestampsEXT(device Device, timestamp_count u32, p_timestamp_infos &CalibratedTimestampInfoKHR, p_timestamps &u64, p_max_deviation &u64) Result

pub type PFN_vkGetCalibratedTimestampsEXT = fn (device Device, timestamp_count u32, p_timestamp_infos &CalibratedTimestampInfoKHR, p_timestamps &u64, p_max_deviation &u64) Result

@[inline]
pub fn get_calibrated_timestamps_ext(device Device,
	timestamp_count u32,
	p_timestamp_infos &CalibratedTimestampInfoKHR,
	p_timestamps &u64,
	p_max_deviation &u64) Result {
	return C.vkGetCalibratedTimestampsEXT(device, timestamp_count, p_timestamp_infos,
		p_timestamps, p_max_deviation)
}

pub const amd_shader_core_properties_spec_version = 2
pub const amd_shader_core_properties_extension_name = c'VK_AMD_shader_core_properties'
// PhysicalDeviceShaderCorePropertiesAMD extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceShaderCorePropertiesAMD = C.VkPhysicalDeviceShaderCorePropertiesAMD

@[typedef]
pub struct C.VkPhysicalDeviceShaderCorePropertiesAMD {
pub mut:
	sType                      StructureType = StructureType.physical_device_shader_core_properties_amd
	pNext                      voidptr       = unsafe { nil }
	shaderEngineCount          u32
	shaderArraysPerEngineCount u32
	computeUnitsPerShaderArray u32
	simdPerComputeUnit         u32
	wavefrontsPerSimd          u32
	wavefrontSize              u32
	sgprsPerSimd               u32
	minSgprAllocation          u32
	maxSgprAllocation          u32
	sgprAllocationGranularity  u32
	vgprsPerSimd               u32
	minVgprAllocation          u32
	maxVgprAllocation          u32
	vgprAllocationGranularity  u32
}

pub const amd_memory_overallocation_behavior_spec_version = 1
pub const amd_memory_overallocation_behavior_extension_name = c'VK_AMD_memory_overallocation_behavior'

pub enum MemoryOverallocationBehaviorAMD as u32 {
	default      = 0
	allowed      = 1
	disallowed   = 2
	max_enum_amd = max_int
}
// DeviceMemoryOverallocationCreateInfoAMD extends VkDeviceCreateInfo
pub type DeviceMemoryOverallocationCreateInfoAMD = C.VkDeviceMemoryOverallocationCreateInfoAMD

@[typedef]
pub struct C.VkDeviceMemoryOverallocationCreateInfoAMD {
pub mut:
	sType                  StructureType = StructureType.device_memory_overallocation_create_info_amd
	pNext                  voidptr       = unsafe { nil }
	overallocationBehavior MemoryOverallocationBehaviorAMD
}

pub const ext_vertex_attribute_divisor_spec_version = 3
pub const ext_vertex_attribute_divisor_extension_name = c'VK_EXT_vertex_attribute_divisor'
// PhysicalDeviceVertexAttributeDivisorPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceVertexAttributeDivisorPropertiesEXT = C.VkPhysicalDeviceVertexAttributeDivisorPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceVertexAttributeDivisorPropertiesEXT {
pub mut:
	sType                  StructureType = StructureType.physical_device_vertex_attribute_divisor_properties_ext
	pNext                  voidptr       = unsafe { nil }
	maxVertexAttribDivisor u32
}

pub type VertexInputBindingDivisorDescriptionEXT = C.VkVertexInputBindingDivisorDescription

pub type PipelineVertexInputDivisorStateCreateInfoEXT = C.VkPipelineVertexInputDivisorStateCreateInfo

pub type PhysicalDeviceVertexAttributeDivisorFeaturesEXT = C.VkPhysicalDeviceVertexAttributeDivisorFeatures

pub const ext_pipeline_creation_feedback_spec_version = 1
pub const ext_pipeline_creation_feedback_extension_name = c'VK_EXT_pipeline_creation_feedback'

pub type PipelineCreationFeedbackFlagBitsEXT = PipelineCreationFeedbackFlagBits

pub type PipelineCreationFeedbackFlagsEXT = u32
pub type PipelineCreationFeedbackCreateInfoEXT = C.VkPipelineCreationFeedbackCreateInfo

pub type PipelineCreationFeedbackEXT = C.VkPipelineCreationFeedback

pub const nv_shader_subgroup_partitioned_spec_version = 1
pub const nv_shader_subgroup_partitioned_extension_name = c'VK_NV_shader_subgroup_partitioned'

pub const nv_compute_shader_derivatives_spec_version = 1
pub const nv_compute_shader_derivatives_extension_name = c'VK_NV_compute_shader_derivatives'

pub type PhysicalDeviceComputeShaderDerivativesFeaturesNV = C.VkPhysicalDeviceComputeShaderDerivativesFeaturesKHR

pub const nv_mesh_shader_spec_version = 1
pub const nv_mesh_shader_extension_name = c'VK_NV_mesh_shader'
// PhysicalDeviceMeshShaderFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMeshShaderFeaturesNV = C.VkPhysicalDeviceMeshShaderFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceMeshShaderFeaturesNV {
pub mut:
	sType      StructureType = StructureType.physical_device_mesh_shader_features_nv
	pNext      voidptr       = unsafe { nil }
	taskShader Bool32
	meshShader Bool32
}

// PhysicalDeviceMeshShaderPropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMeshShaderPropertiesNV = C.VkPhysicalDeviceMeshShaderPropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceMeshShaderPropertiesNV {
pub mut:
	sType                             StructureType = StructureType.physical_device_mesh_shader_properties_nv
	pNext                             voidptr       = unsafe { nil }
	maxDrawMeshTasksCount             u32
	maxTaskWorkGroupInvocations       u32
	maxTaskWorkGroupSize              [3]u32
	maxTaskTotalMemorySize            u32
	maxTaskOutputCount                u32
	maxMeshWorkGroupInvocations       u32
	maxMeshWorkGroupSize              [3]u32
	maxMeshTotalMemorySize            u32
	maxMeshOutputVertices             u32
	maxMeshOutputPrimitives           u32
	maxMeshMultiviewViewCount         u32
	meshOutputPerVertexGranularity    u32
	meshOutputPerPrimitiveGranularity u32
}

pub type DrawMeshTasksIndirectCommandNV = C.VkDrawMeshTasksIndirectCommandNV

@[typedef]
pub struct C.VkDrawMeshTasksIndirectCommandNV {
pub mut:
	taskCount u32
	firstTask u32
}

@[keep_args_alive]
fn C.vkCmdDrawMeshTasksNV(command_buffer CommandBuffer, task_count u32, first_task u32)

pub type PFN_vkCmdDrawMeshTasksNV = fn (command_buffer CommandBuffer, task_count u32, first_task u32)

@[inline]
pub fn cmd_draw_mesh_tasks_nv(command_buffer CommandBuffer,
	task_count u32,
	first_task u32) {
	C.vkCmdDrawMeshTasksNV(command_buffer, task_count, first_task)
}

@[keep_args_alive]
fn C.vkCmdDrawMeshTasksIndirectNV(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, draw_count u32, stride u32)

pub type PFN_vkCmdDrawMeshTasksIndirectNV = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_mesh_tasks_indirect_nv(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	draw_count u32,
	stride u32) {
	C.vkCmdDrawMeshTasksIndirectNV(command_buffer, buffer, offset, draw_count, stride)
}

@[keep_args_alive]
fn C.vkCmdDrawMeshTasksIndirectCountNV(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

pub type PFN_vkCmdDrawMeshTasksIndirectCountNV = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_mesh_tasks_indirect_count_nv(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	count_buffer Buffer,
	count_buffer_offset DeviceSize,
	max_draw_count u32,
	stride u32) {
	C.vkCmdDrawMeshTasksIndirectCountNV(command_buffer, buffer, offset, count_buffer,
		count_buffer_offset, max_draw_count, stride)
}

pub const nv_fragment_shader_barycentric_spec_version = 1
pub const nv_fragment_shader_barycentric_extension_name = c'VK_NV_fragment_shader_barycentric'

pub type PhysicalDeviceFragmentShaderBarycentricFeaturesNV = C.VkPhysicalDeviceFragmentShaderBarycentricFeaturesKHR

pub const nv_shader_image_footprint_spec_version = 2
pub const nv_shader_image_footprint_extension_name = c'VK_NV_shader_image_footprint'
// PhysicalDeviceShaderImageFootprintFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderImageFootprintFeaturesNV = C.VkPhysicalDeviceShaderImageFootprintFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceShaderImageFootprintFeaturesNV {
pub mut:
	sType          StructureType = StructureType.physical_device_shader_image_footprint_features_nv
	pNext          voidptr       = unsafe { nil }
	imageFootprint Bool32
}

pub const nv_scissor_exclusive_spec_version = 2
pub const nv_scissor_exclusive_extension_name = c'VK_NV_scissor_exclusive'
// PipelineViewportExclusiveScissorStateCreateInfoNV extends VkPipelineViewportStateCreateInfo
pub type PipelineViewportExclusiveScissorStateCreateInfoNV = C.VkPipelineViewportExclusiveScissorStateCreateInfoNV

@[typedef]
pub struct C.VkPipelineViewportExclusiveScissorStateCreateInfoNV {
pub mut:
	sType                 StructureType = StructureType.pipeline_viewport_exclusive_scissor_state_create_info_nv
	pNext                 voidptr       = unsafe { nil }
	exclusiveScissorCount u32
	pExclusiveScissors    &Rect2D
}

// PhysicalDeviceExclusiveScissorFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceExclusiveScissorFeaturesNV = C.VkPhysicalDeviceExclusiveScissorFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceExclusiveScissorFeaturesNV {
pub mut:
	sType            StructureType = StructureType.physical_device_exclusive_scissor_features_nv
	pNext            voidptr       = unsafe { nil }
	exclusiveScissor Bool32
}

@[keep_args_alive]
fn C.vkCmdSetExclusiveScissorEnableNV(command_buffer CommandBuffer, first_exclusive_scissor u32, exclusive_scissor_count u32, p_exclusive_scissor_enables &Bool32)

pub type PFN_vkCmdSetExclusiveScissorEnableNV = fn (command_buffer CommandBuffer, first_exclusive_scissor u32, exclusive_scissor_count u32, p_exclusive_scissor_enables &Bool32)

@[inline]
pub fn cmd_set_exclusive_scissor_enable_nv(command_buffer CommandBuffer,
	first_exclusive_scissor u32,
	exclusive_scissor_count u32,
	p_exclusive_scissor_enables &Bool32) {
	C.vkCmdSetExclusiveScissorEnableNV(command_buffer, first_exclusive_scissor, exclusive_scissor_count,
		p_exclusive_scissor_enables)
}

@[keep_args_alive]
fn C.vkCmdSetExclusiveScissorNV(command_buffer CommandBuffer, first_exclusive_scissor u32, exclusive_scissor_count u32, p_exclusive_scissors &Rect2D)

pub type PFN_vkCmdSetExclusiveScissorNV = fn (command_buffer CommandBuffer, first_exclusive_scissor u32, exclusive_scissor_count u32, p_exclusive_scissors &Rect2D)

@[inline]
pub fn cmd_set_exclusive_scissor_nv(command_buffer CommandBuffer,
	first_exclusive_scissor u32,
	exclusive_scissor_count u32,
	p_exclusive_scissors &Rect2D) {
	C.vkCmdSetExclusiveScissorNV(command_buffer, first_exclusive_scissor, exclusive_scissor_count,
		p_exclusive_scissors)
}

pub const nv_device_diagnostic_checkpoints_spec_version = 2
pub const nv_device_diagnostic_checkpoints_extension_name = c'VK_NV_device_diagnostic_checkpoints'
// QueueFamilyCheckpointPropertiesNV extends VkQueueFamilyProperties2
pub type QueueFamilyCheckpointPropertiesNV = C.VkQueueFamilyCheckpointPropertiesNV

@[typedef]
pub struct C.VkQueueFamilyCheckpointPropertiesNV {
pub mut:
	sType                        StructureType = StructureType.queue_family_checkpoint_properties_nv
	pNext                        voidptr       = unsafe { nil }
	checkpointExecutionStageMask PipelineStageFlags
}

pub type CheckpointDataNV = C.VkCheckpointDataNV

@[typedef]
pub struct C.VkCheckpointDataNV {
pub mut:
	sType             StructureType = StructureType.checkpoint_data_nv
	pNext             voidptr       = unsafe { nil }
	stage             PipelineStageFlagBits
	pCheckpointMarker voidptr
}

// QueueFamilyCheckpointProperties2NV extends VkQueueFamilyProperties2
pub type QueueFamilyCheckpointProperties2NV = C.VkQueueFamilyCheckpointProperties2NV

@[typedef]
pub struct C.VkQueueFamilyCheckpointProperties2NV {
pub mut:
	sType                        StructureType = StructureType.queue_family_checkpoint_properties2_nv
	pNext                        voidptr       = unsafe { nil }
	checkpointExecutionStageMask PipelineStageFlags2
}

pub type CheckpointData2NV = C.VkCheckpointData2NV

@[typedef]
pub struct C.VkCheckpointData2NV {
pub mut:
	sType             StructureType = StructureType.checkpoint_data2_nv
	pNext             voidptr       = unsafe { nil }
	stage             PipelineStageFlags2
	pCheckpointMarker voidptr
}

@[keep_args_alive]
fn C.vkCmdSetCheckpointNV(command_buffer CommandBuffer, p_checkpoint_marker voidptr)

pub type PFN_vkCmdSetCheckpointNV = fn (command_buffer CommandBuffer, p_checkpoint_marker voidptr)

@[inline]
pub fn cmd_set_checkpoint_nv(command_buffer CommandBuffer,
	p_checkpoint_marker voidptr) {
	C.vkCmdSetCheckpointNV(command_buffer, p_checkpoint_marker)
}

@[keep_args_alive]
fn C.vkGetQueueCheckpointDataNV(queue Queue, p_checkpoint_data_count &u32, mut p_checkpoint_data CheckpointDataNV)

pub type PFN_vkGetQueueCheckpointDataNV = fn (queue Queue, p_checkpoint_data_count &u32, mut p_checkpoint_data CheckpointDataNV)

@[inline]
pub fn get_queue_checkpoint_data_nv(queue Queue,
	p_checkpoint_data_count &u32,
	mut p_checkpoint_data CheckpointDataNV) {
	C.vkGetQueueCheckpointDataNV(queue, p_checkpoint_data_count, mut p_checkpoint_data)
}

@[keep_args_alive]
fn C.vkGetQueueCheckpointData2NV(queue Queue, p_checkpoint_data_count &u32, mut p_checkpoint_data CheckpointData2NV)

pub type PFN_vkGetQueueCheckpointData2NV = fn (queue Queue, p_checkpoint_data_count &u32, mut p_checkpoint_data CheckpointData2NV)

@[inline]
pub fn get_queue_checkpoint_data2_nv(queue Queue,
	p_checkpoint_data_count &u32,
	mut p_checkpoint_data CheckpointData2NV) {
	C.vkGetQueueCheckpointData2NV(queue, p_checkpoint_data_count, mut p_checkpoint_data)
}

pub const intel_shader_integer_functions_2_spec_version = 1
pub const intel_shader_integer_functions_2_extension_name = c'VK_INTE_shader_integer_functions2'
// PhysicalDeviceShaderIntegerFunctions2FeaturesINTEL extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderIntegerFunctions2FeaturesINTEL = C.VkPhysicalDeviceShaderIntegerFunctions2FeaturesINTEL

@[typedef]
pub struct C.VkPhysicalDeviceShaderIntegerFunctions2FeaturesINTEL {
pub mut:
	sType                   StructureType = StructureType.physical_device_shader_integer_functions2_features_intel
	pNext                   voidptr       = unsafe { nil }
	shaderIntegerFunctions2 Bool32
}

// Pointer to VkPerformanceConfigurationINTEL_T
pub type PerformanceConfigurationINTEL = voidptr

pub const intel_performance_query_spec_version = 2
pub const intel_performance_query_extension_name = c'VK_INTE_performance_query'

pub enum PerformanceConfigurationTypeINTEL as u32 {
	command_queue_metrics_discovery_activated = 0
	max_enum_intel                            = max_int
}

pub enum QueryPoolSamplingModeINTEL as u32 {
	manual         = 0
	max_enum_intel = max_int
}

pub enum PerformanceOverrideTypeINTEL as u32 {
	null_hardware    = 0
	flush_gpu_caches = 1
	max_enum_intel   = max_int
}

pub enum PerformanceParameterTypeINTEL as u32 {
	hw_counters_supported    = 0
	stream_marker_valid_bits = 1
	max_enum_intel           = max_int
}

pub enum PerformanceValueTypeINTEL as u32 {
	uint32         = 0
	uint64         = 1
	float          = 2
	bool           = 3
	string         = 4
	max_enum_intel = max_int
}
pub type PerformanceValueDataINTEL = C.VkPerformanceValueDataINTEL

@[typedef]
pub union C.VkPerformanceValueDataINTEL {
pub mut:
	value32     u32
	value64     u64
	valueFloat  f32
	valueBool   Bool32
	valueString &char
}

pub type PerformanceValueINTEL = C.VkPerformanceValueINTEL

@[typedef]
pub struct C.VkPerformanceValueINTEL {
pub mut:
	type PerformanceValueTypeINTEL
	data PerformanceValueDataINTEL
}

pub type InitializePerformanceApiInfoINTEL = C.VkInitializePerformanceApiInfoINTEL

@[typedef]
pub struct C.VkInitializePerformanceApiInfoINTEL {
pub mut:
	sType     StructureType = StructureType.initialize_performance_api_info_intel
	pNext     voidptr       = unsafe { nil }
	pUserData voidptr       = unsafe { nil }
}

// QueryPoolPerformanceQueryCreateInfoINTEL extends VkQueryPoolCreateInfo
pub type QueryPoolPerformanceQueryCreateInfoINTEL = C.VkQueryPoolPerformanceQueryCreateInfoINTEL

@[typedef]
pub struct C.VkQueryPoolPerformanceQueryCreateInfoINTEL {
pub mut:
	sType                       StructureType = StructureType.query_pool_performance_query_create_info_intel
	pNext                       voidptr       = unsafe { nil }
	performanceCountersSampling QueryPoolSamplingModeINTEL
}

pub type QueryPoolCreateInfoINTEL = C.VkQueryPoolPerformanceQueryCreateInfoINTEL

pub type PerformanceMarkerInfoINTEL = C.VkPerformanceMarkerInfoINTEL

@[typedef]
pub struct C.VkPerformanceMarkerInfoINTEL {
pub mut:
	sType  StructureType = StructureType.performance_marker_info_intel
	pNext  voidptr       = unsafe { nil }
	marker u64
}

pub type PerformanceStreamMarkerInfoINTEL = C.VkPerformanceStreamMarkerInfoINTEL

@[typedef]
pub struct C.VkPerformanceStreamMarkerInfoINTEL {
pub mut:
	sType  StructureType = StructureType.performance_stream_marker_info_intel
	pNext  voidptr       = unsafe { nil }
	marker u32
}

pub type PerformanceOverrideInfoINTEL = C.VkPerformanceOverrideInfoINTEL

@[typedef]
pub struct C.VkPerformanceOverrideInfoINTEL {
pub mut:
	sType     StructureType = StructureType.performance_override_info_intel
	pNext     voidptr       = unsafe { nil }
	type      PerformanceOverrideTypeINTEL
	enable    Bool32
	parameter u64
}

pub type PerformanceConfigurationAcquireInfoINTEL = C.VkPerformanceConfigurationAcquireInfoINTEL

@[typedef]
pub struct C.VkPerformanceConfigurationAcquireInfoINTEL {
pub mut:
	sType StructureType = StructureType.performance_configuration_acquire_info_intel
	pNext voidptr       = unsafe { nil }
	type  PerformanceConfigurationTypeINTEL
}

@[keep_args_alive]
fn C.vkInitializePerformanceApiINTEL(device Device, p_initialize_info &InitializePerformanceApiInfoINTEL) Result

pub type PFN_vkInitializePerformanceApiINTEL = fn (device Device, p_initialize_info &InitializePerformanceApiInfoINTEL) Result

@[inline]
pub fn initialize_performance_api_intel(device Device,
	p_initialize_info &InitializePerformanceApiInfoINTEL) Result {
	return C.vkInitializePerformanceApiINTEL(device, p_initialize_info)
}

@[keep_args_alive]
fn C.vkUninitializePerformanceApiINTEL(device Device)

pub type PFN_vkUninitializePerformanceApiINTEL = fn (device Device)

@[inline]
pub fn uninitialize_performance_api_intel(device Device) {
	C.vkUninitializePerformanceApiINTEL(device)
}

@[keep_args_alive]
fn C.vkCmdSetPerformanceMarkerINTEL(command_buffer CommandBuffer, p_marker_info &PerformanceMarkerInfoINTEL) Result

pub type PFN_vkCmdSetPerformanceMarkerINTEL = fn (command_buffer CommandBuffer, p_marker_info &PerformanceMarkerInfoINTEL) Result

@[inline]
pub fn cmd_set_performance_marker_intel(command_buffer CommandBuffer,
	p_marker_info &PerformanceMarkerInfoINTEL) Result {
	return C.vkCmdSetPerformanceMarkerINTEL(command_buffer, p_marker_info)
}

@[keep_args_alive]
fn C.vkCmdSetPerformanceStreamMarkerINTEL(command_buffer CommandBuffer, p_marker_info &PerformanceStreamMarkerInfoINTEL) Result

pub type PFN_vkCmdSetPerformanceStreamMarkerINTEL = fn (command_buffer CommandBuffer, p_marker_info &PerformanceStreamMarkerInfoINTEL) Result

@[inline]
pub fn cmd_set_performance_stream_marker_intel(command_buffer CommandBuffer,
	p_marker_info &PerformanceStreamMarkerInfoINTEL) Result {
	return C.vkCmdSetPerformanceStreamMarkerINTEL(command_buffer, p_marker_info)
}

@[keep_args_alive]
fn C.vkCmdSetPerformanceOverrideINTEL(command_buffer CommandBuffer, p_override_info &PerformanceOverrideInfoINTEL) Result

pub type PFN_vkCmdSetPerformanceOverrideINTEL = fn (command_buffer CommandBuffer, p_override_info &PerformanceOverrideInfoINTEL) Result

@[inline]
pub fn cmd_set_performance_override_intel(command_buffer CommandBuffer,
	p_override_info &PerformanceOverrideInfoINTEL) Result {
	return C.vkCmdSetPerformanceOverrideINTEL(command_buffer, p_override_info)
}

@[keep_args_alive]
fn C.vkAcquirePerformanceConfigurationINTEL(device Device, p_acquire_info &PerformanceConfigurationAcquireInfoINTEL, p_configuration &PerformanceConfigurationINTEL) Result

pub type PFN_vkAcquirePerformanceConfigurationINTEL = fn (device Device, p_acquire_info &PerformanceConfigurationAcquireInfoINTEL, p_configuration &PerformanceConfigurationINTEL) Result

@[inline]
pub fn acquire_performance_configuration_intel(device Device,
	p_acquire_info &PerformanceConfigurationAcquireInfoINTEL,
	p_configuration &PerformanceConfigurationINTEL) Result {
	return C.vkAcquirePerformanceConfigurationINTEL(device, p_acquire_info, p_configuration)
}

@[keep_args_alive]
fn C.vkReleasePerformanceConfigurationINTEL(device Device, configuration PerformanceConfigurationINTEL) Result

pub type PFN_vkReleasePerformanceConfigurationINTEL = fn (device Device, configuration PerformanceConfigurationINTEL) Result

@[inline]
pub fn release_performance_configuration_intel(device Device,
	configuration PerformanceConfigurationINTEL) Result {
	return C.vkReleasePerformanceConfigurationINTEL(device, configuration)
}

@[keep_args_alive]
fn C.vkQueueSetPerformanceConfigurationINTEL(queue Queue, configuration PerformanceConfigurationINTEL) Result

pub type PFN_vkQueueSetPerformanceConfigurationINTEL = fn (queue Queue, configuration PerformanceConfigurationINTEL) Result

@[inline]
pub fn queue_set_performance_configuration_intel(queue Queue,
	configuration PerformanceConfigurationINTEL) Result {
	return C.vkQueueSetPerformanceConfigurationINTEL(queue, configuration)
}

@[keep_args_alive]
fn C.vkGetPerformanceParameterINTEL(device Device, parameter PerformanceParameterTypeINTEL, mut p_value PerformanceValueINTEL) Result

pub type PFN_vkGetPerformanceParameterINTEL = fn (device Device, parameter PerformanceParameterTypeINTEL, mut p_value PerformanceValueINTEL) Result

@[inline]
pub fn get_performance_parameter_intel(device Device,
	parameter PerformanceParameterTypeINTEL,
	mut p_value PerformanceValueINTEL) Result {
	return C.vkGetPerformanceParameterINTEL(device, parameter, mut p_value)
}

pub const ext_pci_bus_info_spec_version = 2
pub const ext_pci_bus_info_extension_name = c'VK_EXT_pci_bus_info'
// PhysicalDevicePCIBusInfoPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDevicePCIBusInfoPropertiesEXT = C.VkPhysicalDevicePCIBusInfoPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDevicePCIBusInfoPropertiesEXT {
pub mut:
	sType       StructureType = StructureType.physical_device_pci_bus_info_properties_ext
	pNext       voidptr       = unsafe { nil }
	pciDomain   u32
	pciBus      u32
	pciDevice   u32
	pciFunction u32
}

pub const amd_display_native_hdr_spec_version = 1
pub const amd_display_native_hdr_extension_name = c'VK_AMD_display_native_hdr'
// DisplayNativeHdrSurfaceCapabilitiesAMD extends VkSurfaceCapabilities2KHR
pub type DisplayNativeHdrSurfaceCapabilitiesAMD = C.VkDisplayNativeHdrSurfaceCapabilitiesAMD

@[typedef]
pub struct C.VkDisplayNativeHdrSurfaceCapabilitiesAMD {
pub mut:
	sType               StructureType = StructureType.display_native_hdr_surface_capabilities_amd
	pNext               voidptr       = unsafe { nil }
	localDimmingSupport Bool32
}

// SwapchainDisplayNativeHdrCreateInfoAMD extends VkSwapchainCreateInfoKHR
pub type SwapchainDisplayNativeHdrCreateInfoAMD = C.VkSwapchainDisplayNativeHdrCreateInfoAMD

@[typedef]
pub struct C.VkSwapchainDisplayNativeHdrCreateInfoAMD {
pub mut:
	sType              StructureType = StructureType.swapchain_display_native_hdr_create_info_amd
	pNext              voidptr       = unsafe { nil }
	localDimmingEnable Bool32
}

@[keep_args_alive]
fn C.vkSetLocalDimmingAMD(device Device, swap_chain SwapchainKHR, local_dimming_enable Bool32)

pub type PFN_vkSetLocalDimmingAMD = fn (device Device, swap_chain SwapchainKHR, local_dimming_enable Bool32)

@[inline]
pub fn set_local_dimming_amd(device Device,
	swap_chain SwapchainKHR,
	local_dimming_enable Bool32) {
	C.vkSetLocalDimmingAMD(device, swap_chain, local_dimming_enable)
}

pub const ext_fragment_density_map_spec_version = 2
pub const ext_fragment_density_map_extension_name = c'VK_EXT_fragment_density_map'
// PhysicalDeviceFragmentDensityMapFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceFragmentDensityMapFeaturesEXT = C.VkPhysicalDeviceFragmentDensityMapFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceFragmentDensityMapFeaturesEXT {
pub mut:
	sType                                 StructureType = StructureType.physical_device_fragment_density_map_features_ext
	pNext                                 voidptr       = unsafe { nil }
	fragmentDensityMap                    Bool32
	fragmentDensityMapDynamic             Bool32
	fragmentDensityMapNonSubsampledImages Bool32
}

// PhysicalDeviceFragmentDensityMapPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceFragmentDensityMapPropertiesEXT = C.VkPhysicalDeviceFragmentDensityMapPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceFragmentDensityMapPropertiesEXT {
pub mut:
	sType                       StructureType = StructureType.physical_device_fragment_density_map_properties_ext
	pNext                       voidptr       = unsafe { nil }
	minFragmentDensityTexelSize Extent2D
	maxFragmentDensityTexelSize Extent2D
	fragmentDensityInvocations  Bool32
}

// RenderPassFragmentDensityMapCreateInfoEXT extends VkRenderPassCreateInfo,VkRenderPassCreateInfo2
pub type RenderPassFragmentDensityMapCreateInfoEXT = C.VkRenderPassFragmentDensityMapCreateInfoEXT

@[typedef]
pub struct C.VkRenderPassFragmentDensityMapCreateInfoEXT {
pub mut:
	sType                        StructureType = StructureType.render_pass_fragment_density_map_create_info_ext
	pNext                        voidptr       = unsafe { nil }
	fragmentDensityMapAttachment AttachmentReference
}

// RenderingFragmentDensityMapAttachmentInfoEXT extends VkRenderingInfo
pub type RenderingFragmentDensityMapAttachmentInfoEXT = C.VkRenderingFragmentDensityMapAttachmentInfoEXT

@[typedef]
pub struct C.VkRenderingFragmentDensityMapAttachmentInfoEXT {
pub mut:
	sType       StructureType = StructureType.rendering_fragment_density_map_attachment_info_ext
	pNext       voidptr       = unsafe { nil }
	imageView   ImageView
	imageLayout ImageLayout
}

pub const ext_scalar_block_layout_spec_version = 1
pub const ext_scalar_block_layout_extension_name = c'VK_EXT_scalar_block_layout'

pub type PhysicalDeviceScalarBlockLayoutFeaturesEXT = C.VkPhysicalDeviceScalarBlockLayoutFeatures

pub const google_hlsl_functionality_1_spec_version = 1
pub const google_hlsl_functionality_1_extension_name = c'VK_GOOGE_hlsl_functionality1'
// VK_GOOGLE_HLSL_FUNCTIONALITY1_SPEC_VERSION is a deprecated alias
pub const google_hlsl_functionality1_spec_version = google_hlsl_functionality_1_spec_version
// VK_GOOGLE_HLSL_FUNCTIONALITY1_EXTENSION_NAME is a deprecated alias
pub const google_hlsl_functionality1_extension_name = google_hlsl_functionality_1_extension_name

pub const google_decorate_string_spec_version = 1
pub const google_decorate_string_extension_name = c'VK_GOOGE_decorate_string'

pub const ext_subgroup_size_control_spec_version = 2
pub const ext_subgroup_size_control_extension_name = c'VK_EXT_subgroup_size_control'

pub type PhysicalDeviceSubgroupSizeControlFeaturesEXT = C.VkPhysicalDeviceSubgroupSizeControlFeatures

pub type PhysicalDeviceSubgroupSizeControlPropertiesEXT = C.VkPhysicalDeviceSubgroupSizeControlProperties

pub type PipelineShaderStageRequiredSubgroupSizeCreateInfoEXT = C.VkPipelineShaderStageRequiredSubgroupSizeCreateInfo

pub const amd_shader_core_properties_2_spec_version = 1
pub const amd_shader_core_properties_2_extension_name = c'VK_AMD_shader_core_properties2'

pub enum ShaderCorePropertiesFlagBitsAMD as u32 {
	max_enum_amd = max_int
}
pub type ShaderCorePropertiesFlagsAMD = u32

// PhysicalDeviceShaderCoreProperties2AMD extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceShaderCoreProperties2AMD = C.VkPhysicalDeviceShaderCoreProperties2AMD

@[typedef]
pub struct C.VkPhysicalDeviceShaderCoreProperties2AMD {
pub mut:
	sType                  StructureType = StructureType.physical_device_shader_core_properties2_amd
	pNext                  voidptr       = unsafe { nil }
	shaderCoreFeatures     ShaderCorePropertiesFlagsAMD
	activeComputeUnitCount u32
}

pub const amd_device_coherent_memory_spec_version = 1
pub const amd_device_coherent_memory_extension_name = c'VK_AMD_device_coherent_memory'
// PhysicalDeviceCoherentMemoryFeaturesAMD extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCoherentMemoryFeaturesAMD = C.VkPhysicalDeviceCoherentMemoryFeaturesAMD

@[typedef]
pub struct C.VkPhysicalDeviceCoherentMemoryFeaturesAMD {
pub mut:
	sType                StructureType = StructureType.physical_device_coherent_memory_features_amd
	pNext                voidptr       = unsafe { nil }
	deviceCoherentMemory Bool32
}

pub const ext_shader_image_atomic_int64_spec_version = 1
pub const ext_shader_image_atomic_int64_extension_name = c'VK_EXT_shader_image_atomic_int64'
// PhysicalDeviceShaderImageAtomicInt64FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderImageAtomicInt64FeaturesEXT = C.VkPhysicalDeviceShaderImageAtomicInt64FeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderImageAtomicInt64FeaturesEXT {
pub mut:
	sType                   StructureType = StructureType.physical_device_shader_image_atomic_int64_features_ext
	pNext                   voidptr       = unsafe { nil }
	shaderImageInt64Atomics Bool32
	sparseImageInt64Atomics Bool32
}

pub const ext_memory_budget_spec_version = 1
pub const ext_memory_budget_extension_name = c'VK_EXT_memory_budget'
// PhysicalDeviceMemoryBudgetPropertiesEXT extends VkPhysicalDeviceMemoryProperties2
pub type PhysicalDeviceMemoryBudgetPropertiesEXT = C.VkPhysicalDeviceMemoryBudgetPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMemoryBudgetPropertiesEXT {
pub mut:
	sType      StructureType = StructureType.physical_device_memory_budget_properties_ext
	pNext      voidptr       = unsafe { nil }
	heapBudget [max_memory_heaps]DeviceSize
	heapUsage  [max_memory_heaps]DeviceSize
}

pub const ext_memory_priority_spec_version = 1
pub const ext_memory_priority_extension_name = c'VK_EXT_memory_priority'
// PhysicalDeviceMemoryPriorityFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMemoryPriorityFeaturesEXT = C.VkPhysicalDeviceMemoryPriorityFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMemoryPriorityFeaturesEXT {
pub mut:
	sType          StructureType = StructureType.physical_device_memory_priority_features_ext
	pNext          voidptr       = unsafe { nil }
	memoryPriority Bool32
}

// MemoryPriorityAllocateInfoEXT extends VkMemoryAllocateInfo
pub type MemoryPriorityAllocateInfoEXT = C.VkMemoryPriorityAllocateInfoEXT

@[typedef]
pub struct C.VkMemoryPriorityAllocateInfoEXT {
pub mut:
	sType    StructureType = StructureType.memory_priority_allocate_info_ext
	pNext    voidptr       = unsafe { nil }
	priority f32
}

pub const nv_dedicated_allocation_image_aliasing_spec_version = 1
pub const nv_dedicated_allocation_image_aliasing_extension_name = c'VK_NV_dedicated_allocation_image_aliasing'
// PhysicalDeviceDedicatedAllocationImageAliasingFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDedicatedAllocationImageAliasingFeaturesNV = C.VkPhysicalDeviceDedicatedAllocationImageAliasingFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceDedicatedAllocationImageAliasingFeaturesNV {
pub mut:
	sType                            StructureType = StructureType.physical_device_dedicated_allocation_image_aliasing_features_nv
	pNext                            voidptr       = unsafe { nil }
	dedicatedAllocationImageAliasing Bool32
}

pub const ext_buffer_device_address_spec_version = 2
pub const ext_buffer_device_address_extension_name = c'VK_EXT_buffer_device_address'
// PhysicalDeviceBufferDeviceAddressFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceBufferDeviceAddressFeaturesEXT = C.VkPhysicalDeviceBufferDeviceAddressFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceBufferDeviceAddressFeaturesEXT {
pub mut:
	sType                            StructureType = StructureType.physical_device_buffer_device_address_features_ext
	pNext                            voidptr       = unsafe { nil }
	bufferDeviceAddress              Bool32
	bufferDeviceAddressCaptureReplay Bool32
	bufferDeviceAddressMultiDevice   Bool32
}

pub type PhysicalDeviceBufferAddressFeaturesEXT = C.VkPhysicalDeviceBufferDeviceAddressFeaturesEXT

pub type BufferDeviceAddressInfoEXT = C.VkBufferDeviceAddressInfo

// BufferDeviceAddressCreateInfoEXT extends VkBufferCreateInfo
pub type BufferDeviceAddressCreateInfoEXT = C.VkBufferDeviceAddressCreateInfoEXT

@[typedef]
pub struct C.VkBufferDeviceAddressCreateInfoEXT {
pub mut:
	sType         StructureType = StructureType.buffer_device_address_create_info_ext
	pNext         voidptr       = unsafe { nil }
	deviceAddress DeviceAddress
}

@[keep_args_alive]
fn C.vkGetBufferDeviceAddressEXT(device Device, p_info &BufferDeviceAddressInfo) DeviceAddress

pub type PFN_vkGetBufferDeviceAddressEXT = fn (device Device, p_info &BufferDeviceAddressInfo) DeviceAddress

@[inline]
pub fn get_buffer_device_address_ext(device Device,
	p_info &BufferDeviceAddressInfo) DeviceAddress {
	return C.vkGetBufferDeviceAddressEXT(device, p_info)
}

pub const ext_tooling_info_spec_version = 1
pub const ext_tooling_info_extension_name = c'VK_EXT_tooling_info'

pub type ToolPurposeFlagBitsEXT = ToolPurposeFlagBits

pub type ToolPurposeFlagsEXT = u32
pub type PhysicalDeviceToolPropertiesEXT = C.VkPhysicalDeviceToolProperties

@[keep_args_alive]
fn C.vkGetPhysicalDeviceToolPropertiesEXT(physical_device PhysicalDevice, p_tool_count &u32, mut p_tool_properties PhysicalDeviceToolProperties) Result

pub type PFN_vkGetPhysicalDeviceToolPropertiesEXT = fn (physical_device PhysicalDevice, p_tool_count &u32, mut p_tool_properties PhysicalDeviceToolProperties) Result

@[inline]
pub fn get_physical_device_tool_properties_ext(physical_device PhysicalDevice,
	p_tool_count &u32,
	mut p_tool_properties PhysicalDeviceToolProperties) Result {
	return C.vkGetPhysicalDeviceToolPropertiesEXT(physical_device, p_tool_count, mut p_tool_properties)
}

pub const ext_separate_stencil_usage_spec_version = 1
pub const ext_separate_stencil_usage_extension_name = c'VK_EXT_separate_stencil_usage'

pub type ImageStencilUsageCreateInfoEXT = C.VkImageStencilUsageCreateInfo

pub const ext_validation_features_spec_version = 6
pub const ext_validation_features_extension_name = c'VK_EXT_validation_features'

pub enum ValidationFeatureEnableEXT as u32 {
	gpu_assisted                      = 0
	gpu_assisted_reserve_binding_slot = 1
	best_practices                    = 2
	debug_printf                      = 3
	synchronization_validation        = 4
	max_enum_ext                      = max_int
}

pub enum ValidationFeatureDisableEXT as u32 {
	all                     = 0
	shaders                 = 1
	thread_safety           = 2
	api_parameters          = 3
	object_lifetimes        = 4
	core_checks             = 5
	unique_handles          = 6
	shader_validation_cache = 7
	max_enum_ext            = max_int
}
// ValidationFeaturesEXT extends VkInstanceCreateInfo,VkShaderModuleCreateInfo,VkShaderCreateInfoEXT
pub type ValidationFeaturesEXT = C.VkValidationFeaturesEXT

@[typedef]
pub struct C.VkValidationFeaturesEXT {
pub mut:
	sType                          StructureType = StructureType.validation_features_ext
	pNext                          voidptr       = unsafe { nil }
	enabledValidationFeatureCount  u32
	pEnabledValidationFeatures     &ValidationFeatureEnableEXT
	disabledValidationFeatureCount u32
	pDisabledValidationFeatures    &ValidationFeatureDisableEXT
}

pub const nv_cooperative_matrix_spec_version = 1
pub const nv_cooperative_matrix_extension_name = c'VK_NV_cooperative_matrix'

pub type ComponentTypeNV = ComponentTypeKHR

pub type ScopeNV = ScopeKHR

pub type CooperativeMatrixPropertiesNV = C.VkCooperativeMatrixPropertiesNV

@[typedef]
pub struct C.VkCooperativeMatrixPropertiesNV {
pub mut:
	sType StructureType = StructureType.cooperative_matrix_properties_nv
	pNext voidptr       = unsafe { nil }
	MSize u32
	NSize u32
	KSize u32
	AType ComponentTypeNV
	BType ComponentTypeNV
	CType ComponentTypeNV
	DType ComponentTypeNV
	scope ScopeNV
}

// PhysicalDeviceCooperativeMatrixFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCooperativeMatrixFeaturesNV = C.VkPhysicalDeviceCooperativeMatrixFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceCooperativeMatrixFeaturesNV {
pub mut:
	sType                               StructureType = StructureType.physical_device_cooperative_matrix_features_nv
	pNext                               voidptr       = unsafe { nil }
	cooperativeMatrix                   Bool32
	cooperativeMatrixRobustBufferAccess Bool32
}

// PhysicalDeviceCooperativeMatrixPropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceCooperativeMatrixPropertiesNV = C.VkPhysicalDeviceCooperativeMatrixPropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceCooperativeMatrixPropertiesNV {
pub mut:
	sType                            StructureType = StructureType.physical_device_cooperative_matrix_properties_nv
	pNext                            voidptr       = unsafe { nil }
	cooperativeMatrixSupportedStages ShaderStageFlags
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceCooperativeMatrixPropertiesNV(physical_device PhysicalDevice, p_property_count &u32, mut p_properties CooperativeMatrixPropertiesNV) Result

pub type PFN_vkGetPhysicalDeviceCooperativeMatrixPropertiesNV = fn (physical_device PhysicalDevice, p_property_count &u32, mut p_properties CooperativeMatrixPropertiesNV) Result

@[inline]
pub fn get_physical_device_cooperative_matrix_properties_nv(physical_device PhysicalDevice,
	p_property_count &u32,
	mut p_properties CooperativeMatrixPropertiesNV) Result {
	return C.vkGetPhysicalDeviceCooperativeMatrixPropertiesNV(physical_device, p_property_count, mut
		p_properties)
}

pub const nv_coverage_reduction_mode_spec_version = 1
pub const nv_coverage_reduction_mode_extension_name = c'VK_NV_coverage_reduction_mode'

pub enum CoverageReductionModeNV as u32 {
	merge       = 0
	truncate    = 1
	max_enum_nv = max_int
}
pub type PipelineCoverageReductionStateCreateFlagsNV = u32

// PhysicalDeviceCoverageReductionModeFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCoverageReductionModeFeaturesNV = C.VkPhysicalDeviceCoverageReductionModeFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceCoverageReductionModeFeaturesNV {
pub mut:
	sType                 StructureType = StructureType.physical_device_coverage_reduction_mode_features_nv
	pNext                 voidptr       = unsafe { nil }
	coverageReductionMode Bool32
}

// PipelineCoverageReductionStateCreateInfoNV extends VkPipelineMultisampleStateCreateInfo
pub type PipelineCoverageReductionStateCreateInfoNV = C.VkPipelineCoverageReductionStateCreateInfoNV

@[typedef]
pub struct C.VkPipelineCoverageReductionStateCreateInfoNV {
pub mut:
	sType                 StructureType = StructureType.pipeline_coverage_reduction_state_create_info_nv
	pNext                 voidptr       = unsafe { nil }
	flags                 PipelineCoverageReductionStateCreateFlagsNV
	coverageReductionMode CoverageReductionModeNV
}

pub type FramebufferMixedSamplesCombinationNV = C.VkFramebufferMixedSamplesCombinationNV

@[typedef]
pub struct C.VkFramebufferMixedSamplesCombinationNV {
pub mut:
	sType                 StructureType = StructureType.framebuffer_mixed_samples_combination_nv
	pNext                 voidptr       = unsafe { nil }
	coverageReductionMode CoverageReductionModeNV
	rasterizationSamples  SampleCountFlagBits
	depthStencilSamples   SampleCountFlags
	colorSamples          SampleCountFlags
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceSupportedFramebufferMixedSamplesCombinationsNV(physical_device PhysicalDevice, p_combination_count &u32, mut p_combinations FramebufferMixedSamplesCombinationNV) Result

pub type PFN_vkGetPhysicalDeviceSupportedFramebufferMixedSamplesCombinationsNV = fn (physical_device PhysicalDevice, p_combination_count &u32, mut p_combinations FramebufferMixedSamplesCombinationNV) Result

@[inline]
pub fn get_physical_device_supported_framebuffer_mixed_samples_combinations_nv(physical_device PhysicalDevice,
	p_combination_count &u32,
	mut p_combinations FramebufferMixedSamplesCombinationNV) Result {
	return C.vkGetPhysicalDeviceSupportedFramebufferMixedSamplesCombinationsNV(physical_device,
		p_combination_count, mut p_combinations)
}

pub const ext_fragment_shader_interlock_spec_version = 1
pub const ext_fragment_shader_interlock_extension_name = c'VK_EXT_fragment_shader_interlock'
// PhysicalDeviceFragmentShaderInterlockFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceFragmentShaderInterlockFeaturesEXT = C.VkPhysicalDeviceFragmentShaderInterlockFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceFragmentShaderInterlockFeaturesEXT {
pub mut:
	sType                              StructureType = StructureType.physical_device_fragment_shader_interlock_features_ext
	pNext                              voidptr       = unsafe { nil }
	fragmentShaderSampleInterlock      Bool32
	fragmentShaderPixelInterlock       Bool32
	fragmentShaderShadingRateInterlock Bool32
}

pub const ext_ycbcr_image_arrays_spec_version = 1
pub const ext_ycbcr_image_arrays_extension_name = c'VK_EXT_ycbcr_image_arrays'
// PhysicalDeviceYcbcrImageArraysFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceYcbcrImageArraysFeaturesEXT = C.VkPhysicalDeviceYcbcrImageArraysFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceYcbcrImageArraysFeaturesEXT {
pub mut:
	sType            StructureType = StructureType.physical_device_ycbcr_image_arrays_features_ext
	pNext            voidptr       = unsafe { nil }
	ycbcrImageArrays Bool32
}

pub const ext_provoking_vertex_spec_version = 1
pub const ext_provoking_vertex_extension_name = c'VK_EXT_provoking_vertex'

pub enum ProvokingVertexModeEXT as u32 {
	first_vertex = 0
	last_vertex  = 1
	max_enum_ext = max_int
}
// PhysicalDeviceProvokingVertexFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceProvokingVertexFeaturesEXT = C.VkPhysicalDeviceProvokingVertexFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceProvokingVertexFeaturesEXT {
pub mut:
	sType                                     StructureType = StructureType.physical_device_provoking_vertex_features_ext
	pNext                                     voidptr       = unsafe { nil }
	provokingVertexLast                       Bool32
	transformFeedbackPreservesProvokingVertex Bool32
}

// PhysicalDeviceProvokingVertexPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceProvokingVertexPropertiesEXT = C.VkPhysicalDeviceProvokingVertexPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceProvokingVertexPropertiesEXT {
pub mut:
	sType                                                StructureType = StructureType.physical_device_provoking_vertex_properties_ext
	pNext                                                voidptr       = unsafe { nil }
	provokingVertexModePerPipeline                       Bool32
	transformFeedbackPreservesTriangleFanProvokingVertex Bool32
}

// PipelineRasterizationProvokingVertexStateCreateInfoEXT extends VkPipelineRasterizationStateCreateInfo
pub type PipelineRasterizationProvokingVertexStateCreateInfoEXT = C.VkPipelineRasterizationProvokingVertexStateCreateInfoEXT

@[typedef]
pub struct C.VkPipelineRasterizationProvokingVertexStateCreateInfoEXT {
pub mut:
	sType               StructureType = StructureType.pipeline_rasterization_provoking_vertex_state_create_info_ext
	pNext               voidptr       = unsafe { nil }
	provokingVertexMode ProvokingVertexModeEXT
}

pub const ext_headless_surface_spec_version = 1
pub const ext_headless_surface_extension_name = c'VK_EXT_headless_surface'

pub type HeadlessSurfaceCreateFlagsEXT = u32
pub type HeadlessSurfaceCreateInfoEXT = C.VkHeadlessSurfaceCreateInfoEXT

@[typedef]
pub struct C.VkHeadlessSurfaceCreateInfoEXT {
pub mut:
	sType StructureType = StructureType.headless_surface_create_info_ext
	pNext voidptr       = unsafe { nil }
	flags HeadlessSurfaceCreateFlagsEXT
}

@[keep_args_alive]
fn C.vkCreateHeadlessSurfaceEXT(instance Instance, p_create_info &HeadlessSurfaceCreateInfoEXT, p_allocator &AllocationCallbacks, p_surface &SurfaceKHR) Result

pub type PFN_vkCreateHeadlessSurfaceEXT = fn (instance Instance, p_create_info &HeadlessSurfaceCreateInfoEXT, p_allocator &AllocationCallbacks, p_surface &SurfaceKHR) Result

@[inline]
pub fn create_headless_surface_ext(instance Instance,
	p_create_info &HeadlessSurfaceCreateInfoEXT,
	p_allocator &AllocationCallbacks,
	p_surface &SurfaceKHR) Result {
	return C.vkCreateHeadlessSurfaceEXT(instance, p_create_info, p_allocator, p_surface)
}

pub const ext_line_rasterization_spec_version = 1
pub const ext_line_rasterization_extension_name = c'VK_EXT_line_rasterization'

pub type LineRasterizationModeEXT = LineRasterizationMode

pub type PhysicalDeviceLineRasterizationFeaturesEXT = C.VkPhysicalDeviceLineRasterizationFeatures

pub type PhysicalDeviceLineRasterizationPropertiesEXT = C.VkPhysicalDeviceLineRasterizationProperties

pub type PipelineRasterizationLineStateCreateInfoEXT = C.VkPipelineRasterizationLineStateCreateInfo

@[keep_args_alive]
fn C.vkCmdSetLineStippleEXT(command_buffer CommandBuffer, line_stipple_factor u32, line_stipple_pattern u16)

pub type PFN_vkCmdSetLineStippleEXT = fn (command_buffer CommandBuffer, line_stipple_factor u32, line_stipple_pattern u16)

@[inline]
pub fn cmd_set_line_stipple_ext(command_buffer CommandBuffer,
	line_stipple_factor u32,
	line_stipple_pattern u16) {
	C.vkCmdSetLineStippleEXT(command_buffer, line_stipple_factor, line_stipple_pattern)
}

pub const ext_shader_atomic_float_spec_version = 1
pub const ext_shader_atomic_float_extension_name = c'VK_EXT_shader_atomic_float'
// PhysicalDeviceShaderAtomicFloatFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderAtomicFloatFeaturesEXT = C.VkPhysicalDeviceShaderAtomicFloatFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderAtomicFloatFeaturesEXT {
pub mut:
	sType                        StructureType = StructureType.physical_device_shader_atomic_float_features_ext
	pNext                        voidptr       = unsafe { nil }
	shaderBufferFloat32Atomics   Bool32
	shaderBufferFloat32AtomicAdd Bool32
	shaderBufferFloat64Atomics   Bool32
	shaderBufferFloat64AtomicAdd Bool32
	shaderSharedFloat32Atomics   Bool32
	shaderSharedFloat32AtomicAdd Bool32
	shaderSharedFloat64Atomics   Bool32
	shaderSharedFloat64AtomicAdd Bool32
	shaderImageFloat32Atomics    Bool32
	shaderImageFloat32AtomicAdd  Bool32
	sparseImageFloat32Atomics    Bool32
	sparseImageFloat32AtomicAdd  Bool32
}

pub const ext_host_query_reset_spec_version = 1
pub const ext_host_query_reset_extension_name = c'VK_EXT_host_query_reset'

pub type PhysicalDeviceHostQueryResetFeaturesEXT = C.VkPhysicalDeviceHostQueryResetFeatures

@[keep_args_alive]
fn C.vkResetQueryPoolEXT(device Device, query_pool QueryPool, first_query u32, query_count u32)

pub type PFN_vkResetQueryPoolEXT = fn (device Device, query_pool QueryPool, first_query u32, query_count u32)

@[inline]
pub fn reset_query_pool_ext(device Device,
	query_pool QueryPool,
	first_query u32,
	query_count u32) {
	C.vkResetQueryPoolEXT(device, query_pool, first_query, query_count)
}

pub const ext_index_type_uint8_spec_version = 1
pub const ext_index_type_uint8_extension_name = c'VK_EXT_index_type_uint8'

pub type PhysicalDeviceIndexTypeUint8FeaturesEXT = C.VkPhysicalDeviceIndexTypeUint8Features

pub const ext_extended_dynamic_state_spec_version = 1
pub const ext_extended_dynamic_state_extension_name = c'VK_EXT_extended_dynamic_state'
// PhysicalDeviceExtendedDynamicStateFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceExtendedDynamicStateFeaturesEXT = C.VkPhysicalDeviceExtendedDynamicStateFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceExtendedDynamicStateFeaturesEXT {
pub mut:
	sType                StructureType = StructureType.physical_device_extended_dynamic_state_features_ext
	pNext                voidptr       = unsafe { nil }
	extendedDynamicState Bool32
}

@[keep_args_alive]
fn C.vkCmdSetCullModeEXT(command_buffer CommandBuffer, cull_mode CullModeFlags)

pub type PFN_vkCmdSetCullModeEXT = fn (command_buffer CommandBuffer, cull_mode CullModeFlags)

@[inline]
pub fn cmd_set_cull_mode_ext(command_buffer CommandBuffer,
	cull_mode CullModeFlags) {
	C.vkCmdSetCullModeEXT(command_buffer, cull_mode)
}

@[keep_args_alive]
fn C.vkCmdSetFrontFaceEXT(command_buffer CommandBuffer, front_face FrontFace)

pub type PFN_vkCmdSetFrontFaceEXT = fn (command_buffer CommandBuffer, front_face FrontFace)

@[inline]
pub fn cmd_set_front_face_ext(command_buffer CommandBuffer,
	front_face FrontFace) {
	C.vkCmdSetFrontFaceEXT(command_buffer, front_face)
}

@[keep_args_alive]
fn C.vkCmdSetPrimitiveTopologyEXT(command_buffer CommandBuffer, primitive_topology PrimitiveTopology)

pub type PFN_vkCmdSetPrimitiveTopologyEXT = fn (command_buffer CommandBuffer, primitive_topology PrimitiveTopology)

@[inline]
pub fn cmd_set_primitive_topology_ext(command_buffer CommandBuffer,
	primitive_topology PrimitiveTopology) {
	C.vkCmdSetPrimitiveTopologyEXT(command_buffer, primitive_topology)
}

@[keep_args_alive]
fn C.vkCmdSetViewportWithCountEXT(command_buffer CommandBuffer, viewport_count u32, p_viewports &Viewport)

pub type PFN_vkCmdSetViewportWithCountEXT = fn (command_buffer CommandBuffer, viewport_count u32, p_viewports &Viewport)

@[inline]
pub fn cmd_set_viewport_with_count_ext(command_buffer CommandBuffer,
	viewport_count u32,
	p_viewports &Viewport) {
	C.vkCmdSetViewportWithCountEXT(command_buffer, viewport_count, p_viewports)
}

@[keep_args_alive]
fn C.vkCmdSetScissorWithCountEXT(command_buffer CommandBuffer, scissor_count u32, p_scissors &Rect2D)

pub type PFN_vkCmdSetScissorWithCountEXT = fn (command_buffer CommandBuffer, scissor_count u32, p_scissors &Rect2D)

@[inline]
pub fn cmd_set_scissor_with_count_ext(command_buffer CommandBuffer,
	scissor_count u32,
	p_scissors &Rect2D) {
	C.vkCmdSetScissorWithCountEXT(command_buffer, scissor_count, p_scissors)
}

@[keep_args_alive]
fn C.vkCmdBindVertexBuffers2EXT(command_buffer CommandBuffer, first_binding u32, binding_count u32, p_buffers &Buffer, p_offsets &DeviceSize, p_sizes &DeviceSize, p_strides &DeviceSize)

pub type PFN_vkCmdBindVertexBuffers2EXT = fn (command_buffer CommandBuffer, first_binding u32, binding_count u32, p_buffers &Buffer, p_offsets &DeviceSize, p_sizes &DeviceSize, p_strides &DeviceSize)

@[inline]
pub fn cmd_bind_vertex_buffers2_ext(command_buffer CommandBuffer,
	first_binding u32,
	binding_count u32,
	p_buffers &Buffer,
	p_offsets &DeviceSize,
	p_sizes &DeviceSize,
	p_strides &DeviceSize) {
	C.vkCmdBindVertexBuffers2EXT(command_buffer, first_binding, binding_count, p_buffers,
		p_offsets, p_sizes, p_strides)
}

@[keep_args_alive]
fn C.vkCmdSetDepthTestEnableEXT(command_buffer CommandBuffer, depth_test_enable Bool32)

pub type PFN_vkCmdSetDepthTestEnableEXT = fn (command_buffer CommandBuffer, depth_test_enable Bool32)

@[inline]
pub fn cmd_set_depth_test_enable_ext(command_buffer CommandBuffer,
	depth_test_enable Bool32) {
	C.vkCmdSetDepthTestEnableEXT(command_buffer, depth_test_enable)
}

@[keep_args_alive]
fn C.vkCmdSetDepthWriteEnableEXT(command_buffer CommandBuffer, depth_write_enable Bool32)

pub type PFN_vkCmdSetDepthWriteEnableEXT = fn (command_buffer CommandBuffer, depth_write_enable Bool32)

@[inline]
pub fn cmd_set_depth_write_enable_ext(command_buffer CommandBuffer,
	depth_write_enable Bool32) {
	C.vkCmdSetDepthWriteEnableEXT(command_buffer, depth_write_enable)
}

@[keep_args_alive]
fn C.vkCmdSetDepthCompareOpEXT(command_buffer CommandBuffer, depth_compare_op CompareOp)

pub type PFN_vkCmdSetDepthCompareOpEXT = fn (command_buffer CommandBuffer, depth_compare_op CompareOp)

@[inline]
pub fn cmd_set_depth_compare_op_ext(command_buffer CommandBuffer,
	depth_compare_op CompareOp) {
	C.vkCmdSetDepthCompareOpEXT(command_buffer, depth_compare_op)
}

@[keep_args_alive]
fn C.vkCmdSetDepthBoundsTestEnableEXT(command_buffer CommandBuffer, depth_bounds_test_enable Bool32)

pub type PFN_vkCmdSetDepthBoundsTestEnableEXT = fn (command_buffer CommandBuffer, depth_bounds_test_enable Bool32)

@[inline]
pub fn cmd_set_depth_bounds_test_enable_ext(command_buffer CommandBuffer,
	depth_bounds_test_enable Bool32) {
	C.vkCmdSetDepthBoundsTestEnableEXT(command_buffer, depth_bounds_test_enable)
}

@[keep_args_alive]
fn C.vkCmdSetStencilTestEnableEXT(command_buffer CommandBuffer, stencil_test_enable Bool32)

pub type PFN_vkCmdSetStencilTestEnableEXT = fn (command_buffer CommandBuffer, stencil_test_enable Bool32)

@[inline]
pub fn cmd_set_stencil_test_enable_ext(command_buffer CommandBuffer,
	stencil_test_enable Bool32) {
	C.vkCmdSetStencilTestEnableEXT(command_buffer, stencil_test_enable)
}

@[keep_args_alive]
fn C.vkCmdSetStencilOpEXT(command_buffer CommandBuffer, face_mask StencilFaceFlags, fail_op StencilOp, pass_op StencilOp, depth_fail_op StencilOp, compare_op CompareOp)

pub type PFN_vkCmdSetStencilOpEXT = fn (command_buffer CommandBuffer, face_mask StencilFaceFlags, fail_op StencilOp, pass_op StencilOp, depth_fail_op StencilOp, compare_op CompareOp)

@[inline]
pub fn cmd_set_stencil_op_ext(command_buffer CommandBuffer,
	face_mask StencilFaceFlags,
	fail_op StencilOp,
	pass_op StencilOp,
	depth_fail_op StencilOp,
	compare_op CompareOp) {
	C.vkCmdSetStencilOpEXT(command_buffer, face_mask, fail_op, pass_op, depth_fail_op,
		compare_op)
}

pub const ext_host_image_copy_spec_version = 1
pub const ext_host_image_copy_extension_name = c'VK_EXT_host_image_copy'

pub type HostImageCopyFlagBitsEXT = HostImageCopyFlagBits

pub type HostImageCopyFlagsEXT = u32
pub type PhysicalDeviceHostImageCopyFeaturesEXT = C.VkPhysicalDeviceHostImageCopyFeatures

pub type PhysicalDeviceHostImageCopyPropertiesEXT = C.VkPhysicalDeviceHostImageCopyProperties

pub type MemoryToImageCopyEXT = C.VkMemoryToImageCopy

pub type ImageToMemoryCopyEXT = C.VkImageToMemoryCopy

pub type CopyMemoryToImageInfoEXT = C.VkCopyMemoryToImageInfo

pub type CopyImageToMemoryInfoEXT = C.VkCopyImageToMemoryInfo

pub type CopyImageToImageInfoEXT = C.VkCopyImageToImageInfo

pub type HostImageLayoutTransitionInfoEXT = C.VkHostImageLayoutTransitionInfo

pub type SubresourceHostMemcpySizeEXT = C.VkSubresourceHostMemcpySize

pub type HostImageCopyDevicePerformanceQueryEXT = C.VkHostImageCopyDevicePerformanceQuery

pub type SubresourceLayout2EXT = C.VkSubresourceLayout2

pub type ImageSubresource2EXT = C.VkImageSubresource2

@[keep_args_alive]
fn C.vkCopyMemoryToImageEXT(device Device, p_copy_memory_to_image_info &CopyMemoryToImageInfo) Result

pub type PFN_vkCopyMemoryToImageEXT = fn (device Device, p_copy_memory_to_image_info &CopyMemoryToImageInfo) Result

@[inline]
pub fn copy_memory_to_image_ext(device Device,
	p_copy_memory_to_image_info &CopyMemoryToImageInfo) Result {
	return C.vkCopyMemoryToImageEXT(device, p_copy_memory_to_image_info)
}

@[keep_args_alive]
fn C.vkCopyImageToMemoryEXT(device Device, p_copy_image_to_memory_info &CopyImageToMemoryInfo) Result

pub type PFN_vkCopyImageToMemoryEXT = fn (device Device, p_copy_image_to_memory_info &CopyImageToMemoryInfo) Result

@[inline]
pub fn copy_image_to_memory_ext(device Device,
	p_copy_image_to_memory_info &CopyImageToMemoryInfo) Result {
	return C.vkCopyImageToMemoryEXT(device, p_copy_image_to_memory_info)
}

@[keep_args_alive]
fn C.vkCopyImageToImageEXT(device Device, p_copy_image_to_image_info &CopyImageToImageInfo) Result

pub type PFN_vkCopyImageToImageEXT = fn (device Device, p_copy_image_to_image_info &CopyImageToImageInfo) Result

@[inline]
pub fn copy_image_to_image_ext(device Device,
	p_copy_image_to_image_info &CopyImageToImageInfo) Result {
	return C.vkCopyImageToImageEXT(device, p_copy_image_to_image_info)
}

@[keep_args_alive]
fn C.vkTransitionImageLayoutEXT(device Device, transition_count u32, p_transitions &HostImageLayoutTransitionInfo) Result

pub type PFN_vkTransitionImageLayoutEXT = fn (device Device, transition_count u32, p_transitions &HostImageLayoutTransitionInfo) Result

@[inline]
pub fn transition_image_layout_ext(device Device,
	transition_count u32,
	p_transitions &HostImageLayoutTransitionInfo) Result {
	return C.vkTransitionImageLayoutEXT(device, transition_count, p_transitions)
}

@[keep_args_alive]
fn C.vkGetImageSubresourceLayout2EXT(device Device, image Image, p_subresource &ImageSubresource2, mut p_layout SubresourceLayout2)

pub type PFN_vkGetImageSubresourceLayout2EXT = fn (device Device, image Image, p_subresource &ImageSubresource2, mut p_layout SubresourceLayout2)

@[inline]
pub fn get_image_subresource_layout2_ext(device Device,
	image Image,
	p_subresource &ImageSubresource2,
	mut p_layout SubresourceLayout2) {
	C.vkGetImageSubresourceLayout2EXT(device, image, p_subresource, mut p_layout)
}

pub const ext_map_memory_placed_spec_version = 1
pub const ext_map_memory_placed_extension_name = c'VK_EXT_map_memory_placed'
// PhysicalDeviceMapMemoryPlacedFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMapMemoryPlacedFeaturesEXT = C.VkPhysicalDeviceMapMemoryPlacedFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMapMemoryPlacedFeaturesEXT {
pub mut:
	sType                StructureType = StructureType.physical_device_map_memory_placed_features_ext
	pNext                voidptr       = unsafe { nil }
	memoryMapPlaced      Bool32
	memoryMapRangePlaced Bool32
	memoryUnmapReserve   Bool32
}

// PhysicalDeviceMapMemoryPlacedPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMapMemoryPlacedPropertiesEXT = C.VkPhysicalDeviceMapMemoryPlacedPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMapMemoryPlacedPropertiesEXT {
pub mut:
	sType                       StructureType = StructureType.physical_device_map_memory_placed_properties_ext
	pNext                       voidptr       = unsafe { nil }
	minPlacedMemoryMapAlignment DeviceSize
}

// MemoryMapPlacedInfoEXT extends VkMemoryMapInfo
pub type MemoryMapPlacedInfoEXT = C.VkMemoryMapPlacedInfoEXT

@[typedef]
pub struct C.VkMemoryMapPlacedInfoEXT {
pub mut:
	sType          StructureType = StructureType.memory_map_placed_info_ext
	pNext          voidptr       = unsafe { nil }
	pPlacedAddress voidptr
}

pub const ext_shader_atomic_float_2_spec_version = 1
pub const ext_shader_atomic_float_2_extension_name = c'VK_EXT_shader_atomic_float2'
// PhysicalDeviceShaderAtomicFloat2FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderAtomicFloat2FeaturesEXT = C.VkPhysicalDeviceShaderAtomicFloat2FeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderAtomicFloat2FeaturesEXT {
pub mut:
	sType                           StructureType = StructureType.physical_device_shader_atomic_float2_features_ext
	pNext                           voidptr       = unsafe { nil }
	shaderBufferFloat16Atomics      Bool32
	shaderBufferFloat16AtomicAdd    Bool32
	shaderBufferFloat16AtomicMinMax Bool32
	shaderBufferFloat32AtomicMinMax Bool32
	shaderBufferFloat64AtomicMinMax Bool32
	shaderSharedFloat16Atomics      Bool32
	shaderSharedFloat16AtomicAdd    Bool32
	shaderSharedFloat16AtomicMinMax Bool32
	shaderSharedFloat32AtomicMinMax Bool32
	shaderSharedFloat64AtomicMinMax Bool32
	shaderImageFloat32AtomicMinMax  Bool32
	sparseImageFloat32AtomicMinMax  Bool32
}

pub const ext_surface_maintenance_1_spec_version = 1
pub const ext_surface_maintenance_1_extension_name = c'VK_EXT_surface_maintenance1'

pub type PresentScalingFlagBitsEXT = PresentScalingFlagBitsKHR

pub type PresentScalingFlagsEXT = u32
pub type PresentGravityFlagBitsEXT = PresentGravityFlagBitsKHR

pub type PresentGravityFlagsEXT = u32
pub type SurfacePresentModeEXT = C.VkSurfacePresentModeKHR

pub type SurfacePresentScalingCapabilitiesEXT = C.VkSurfacePresentScalingCapabilitiesKHR

pub type SurfacePresentModeCompatibilityEXT = C.VkSurfacePresentModeCompatibilityKHR

pub const ext_swapchain_maintenance_1_spec_version = 1
pub const ext_swapchain_maintenance_1_extension_name = c'VK_EXT_swapchain_maintenance1'

pub type PhysicalDeviceSwapchainMaintenance1FeaturesEXT = C.VkPhysicalDeviceSwapchainMaintenance1FeaturesKHR

pub type SwapchainPresentFenceInfoEXT = C.VkSwapchainPresentFenceInfoKHR

pub type SwapchainPresentModesCreateInfoEXT = C.VkSwapchainPresentModesCreateInfoKHR

pub type SwapchainPresentModeInfoEXT = C.VkSwapchainPresentModeInfoKHR

pub type SwapchainPresentScalingCreateInfoEXT = C.VkSwapchainPresentScalingCreateInfoKHR

pub type ReleaseSwapchainImagesInfoEXT = C.VkReleaseSwapchainImagesInfoKHR

@[keep_args_alive]
fn C.vkReleaseSwapchainImagesEXT(device Device, p_release_info &ReleaseSwapchainImagesInfoKHR) Result

pub type PFN_vkReleaseSwapchainImagesEXT = fn (device Device, p_release_info &ReleaseSwapchainImagesInfoKHR) Result

@[inline]
pub fn release_swapchain_images_ext(device Device,
	p_release_info &ReleaseSwapchainImagesInfoKHR) Result {
	return C.vkReleaseSwapchainImagesEXT(device, p_release_info)
}

pub const ext_shader_demote_to_helper_invocation_spec_version = 1
pub const ext_shader_demote_to_helper_invocation_extension_name = c'VK_EXT_shader_demote_to_helper_invocation'

pub type PhysicalDeviceShaderDemoteToHelperInvocationFeaturesEXT = C.VkPhysicalDeviceShaderDemoteToHelperInvocationFeatures

// Pointer to VkIndirectCommandsLayoutNV_T
pub type IndirectCommandsLayoutNV = voidptr

pub const nv_device_generated_commands_spec_version = 3
pub const nv_device_generated_commands_extension_name = c'VK_NV_device_generated_commands'

pub enum IndirectCommandsTokenTypeNV as u32 {
	shader_group    = 0
	state_flags     = 1
	index_buffer    = 2
	vertex_buffer   = 3
	push_constant   = 4
	draw_indexed    = 5
	draw            = 6
	draw_tasks      = 7
	draw_mesh_tasks = 1000328000
	pipeline        = 1000428003
	dispatch        = 1000428004
	max_enum_nv     = max_int
}

pub enum IndirectStateFlagBitsNV as u32 {
	frontface   = u32(0x00000001)
	max_enum_nv = max_int
}
pub type IndirectStateFlagsNV = u32

pub enum IndirectCommandsLayoutUsageFlagBitsNV as u32 {
	explicit_preprocess = u32(0x00000001)
	indexed_sequences   = u32(0x00000002)
	unordered_sequences = u32(0x00000004)
	max_enum_nv         = max_int
}
pub type IndirectCommandsLayoutUsageFlagsNV = u32

// PhysicalDeviceDeviceGeneratedCommandsPropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceDeviceGeneratedCommandsPropertiesNV = C.VkPhysicalDeviceDeviceGeneratedCommandsPropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceDeviceGeneratedCommandsPropertiesNV {
pub mut:
	sType                                    StructureType = StructureType.physical_device_device_generated_commands_properties_nv
	pNext                                    voidptr       = unsafe { nil }
	maxGraphicsShaderGroupCount              u32
	maxIndirectSequenceCount                 u32
	maxIndirectCommandsTokenCount            u32
	maxIndirectCommandsStreamCount           u32
	maxIndirectCommandsTokenOffset           u32
	maxIndirectCommandsStreamStride          u32
	minSequencesCountBufferOffsetAlignment   u32
	minSequencesIndexBufferOffsetAlignment   u32
	minIndirectCommandsBufferOffsetAlignment u32
}

// PhysicalDeviceDeviceGeneratedCommandsFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDeviceGeneratedCommandsFeaturesNV = C.VkPhysicalDeviceDeviceGeneratedCommandsFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceDeviceGeneratedCommandsFeaturesNV {
pub mut:
	sType                   StructureType = StructureType.physical_device_device_generated_commands_features_nv
	pNext                   voidptr       = unsafe { nil }
	deviceGeneratedCommands Bool32
}

pub type GraphicsShaderGroupCreateInfoNV = C.VkGraphicsShaderGroupCreateInfoNV

@[typedef]
pub struct C.VkGraphicsShaderGroupCreateInfoNV {
pub mut:
	sType              StructureType = StructureType.graphics_shader_group_create_info_nv
	pNext              voidptr       = unsafe { nil }
	stageCount         u32
	pStages            &PipelineShaderStageCreateInfo
	pVertexInputState  &PipelineVertexInputStateCreateInfo
	pTessellationState &PipelineTessellationStateCreateInfo
}

// GraphicsPipelineShaderGroupsCreateInfoNV extends VkGraphicsPipelineCreateInfo
pub type GraphicsPipelineShaderGroupsCreateInfoNV = C.VkGraphicsPipelineShaderGroupsCreateInfoNV

@[typedef]
pub struct C.VkGraphicsPipelineShaderGroupsCreateInfoNV {
pub mut:
	sType         StructureType = StructureType.graphics_pipeline_shader_groups_create_info_nv
	pNext         voidptr       = unsafe { nil }
	groupCount    u32
	pGroups       &GraphicsShaderGroupCreateInfoNV
	pipelineCount u32
	pPipelines    &Pipeline
}

pub type BindShaderGroupIndirectCommandNV = C.VkBindShaderGroupIndirectCommandNV

@[typedef]
pub struct C.VkBindShaderGroupIndirectCommandNV {
pub mut:
	groupIndex u32
}

pub type BindIndexBufferIndirectCommandNV = C.VkBindIndexBufferIndirectCommandNV

@[typedef]
pub struct C.VkBindIndexBufferIndirectCommandNV {
pub mut:
	bufferAddress DeviceAddress
	size          u32
	indexType     IndexType
}

pub type BindVertexBufferIndirectCommandNV = C.VkBindVertexBufferIndirectCommandNV

@[typedef]
pub struct C.VkBindVertexBufferIndirectCommandNV {
pub mut:
	bufferAddress DeviceAddress
	size          u32
	stride        u32
}

pub type SetStateFlagsIndirectCommandNV = C.VkSetStateFlagsIndirectCommandNV

@[typedef]
pub struct C.VkSetStateFlagsIndirectCommandNV {
pub mut:
	data u32
}

pub type IndirectCommandsStreamNV = C.VkIndirectCommandsStreamNV

@[typedef]
pub struct C.VkIndirectCommandsStreamNV {
pub mut:
	buffer Buffer
	offset DeviceSize
}

pub type IndirectCommandsLayoutTokenNV = C.VkIndirectCommandsLayoutTokenNV

@[typedef]
pub struct C.VkIndirectCommandsLayoutTokenNV {
pub mut:
	sType                        StructureType = StructureType.indirect_commands_layout_token_nv
	pNext                        voidptr       = unsafe { nil }
	tokenType                    IndirectCommandsTokenTypeNV
	stream                       u32
	offset                       u32
	vertexBindingUnit            u32
	vertexDynamicStride          Bool32
	pushconstantPipelineLayout   PipelineLayout
	pushconstantShaderStageFlags ShaderStageFlags
	pushconstantOffset           u32
	pushconstantSize             u32
	indirectStateFlags           IndirectStateFlagsNV
	indexTypeCount               u32
	pIndexTypes                  &IndexType
	pIndexTypeValues             &u32
}

pub type IndirectCommandsLayoutCreateInfoNV = C.VkIndirectCommandsLayoutCreateInfoNV

@[typedef]
pub struct C.VkIndirectCommandsLayoutCreateInfoNV {
pub mut:
	sType             StructureType = StructureType.indirect_commands_layout_create_info_nv
	pNext             voidptr       = unsafe { nil }
	flags             IndirectCommandsLayoutUsageFlagsNV
	pipelineBindPoint PipelineBindPoint
	tokenCount        u32
	pTokens           &IndirectCommandsLayoutTokenNV
	streamCount       u32
	pStreamStrides    &u32
}

pub type GeneratedCommandsInfoNV = C.VkGeneratedCommandsInfoNV

@[typedef]
pub struct C.VkGeneratedCommandsInfoNV {
pub mut:
	sType                  StructureType = StructureType.generated_commands_info_nv
	pNext                  voidptr       = unsafe { nil }
	pipelineBindPoint      PipelineBindPoint
	pipeline               Pipeline
	indirectCommandsLayout IndirectCommandsLayoutNV
	streamCount            u32
	pStreams               &IndirectCommandsStreamNV
	sequencesCount         u32
	preprocessBuffer       Buffer
	preprocessOffset       DeviceSize
	preprocessSize         DeviceSize
	sequencesCountBuffer   Buffer
	sequencesCountOffset   DeviceSize
	sequencesIndexBuffer   Buffer
	sequencesIndexOffset   DeviceSize
}

pub type GeneratedCommandsMemoryRequirementsInfoNV = C.VkGeneratedCommandsMemoryRequirementsInfoNV

@[typedef]
pub struct C.VkGeneratedCommandsMemoryRequirementsInfoNV {
pub mut:
	sType                  StructureType = StructureType.generated_commands_memory_requirements_info_nv
	pNext                  voidptr       = unsafe { nil }
	pipelineBindPoint      PipelineBindPoint
	pipeline               Pipeline
	indirectCommandsLayout IndirectCommandsLayoutNV
	maxSequencesCount      u32
}

@[keep_args_alive]
fn C.vkGetGeneratedCommandsMemoryRequirementsNV(device Device, p_info &GeneratedCommandsMemoryRequirementsInfoNV, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetGeneratedCommandsMemoryRequirementsNV = fn (device Device, p_info &GeneratedCommandsMemoryRequirementsInfoNV, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_generated_commands_memory_requirements_nv(device Device,
	p_info &GeneratedCommandsMemoryRequirementsInfoNV,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetGeneratedCommandsMemoryRequirementsNV(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkCmdPreprocessGeneratedCommandsNV(command_buffer CommandBuffer, p_generated_commands_info &GeneratedCommandsInfoNV)

pub type PFN_vkCmdPreprocessGeneratedCommandsNV = fn (command_buffer CommandBuffer, p_generated_commands_info &GeneratedCommandsInfoNV)

@[inline]
pub fn cmd_preprocess_generated_commands_nv(command_buffer CommandBuffer,
	p_generated_commands_info &GeneratedCommandsInfoNV) {
	C.vkCmdPreprocessGeneratedCommandsNV(command_buffer, p_generated_commands_info)
}

@[keep_args_alive]
fn C.vkCmdExecuteGeneratedCommandsNV(command_buffer CommandBuffer, is_preprocessed Bool32, p_generated_commands_info &GeneratedCommandsInfoNV)

pub type PFN_vkCmdExecuteGeneratedCommandsNV = fn (command_buffer CommandBuffer, is_preprocessed Bool32, p_generated_commands_info &GeneratedCommandsInfoNV)

@[inline]
pub fn cmd_execute_generated_commands_nv(command_buffer CommandBuffer,
	is_preprocessed Bool32,
	p_generated_commands_info &GeneratedCommandsInfoNV) {
	C.vkCmdExecuteGeneratedCommandsNV(command_buffer, is_preprocessed, p_generated_commands_info)
}

@[keep_args_alive]
fn C.vkCmdBindPipelineShaderGroupNV(command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, pipeline Pipeline, group_index u32)

pub type PFN_vkCmdBindPipelineShaderGroupNV = fn (command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, pipeline Pipeline, group_index u32)

@[inline]
pub fn cmd_bind_pipeline_shader_group_nv(command_buffer CommandBuffer,
	pipeline_bind_point PipelineBindPoint,
	pipeline Pipeline,
	group_index u32) {
	C.vkCmdBindPipelineShaderGroupNV(command_buffer, pipeline_bind_point, pipeline, group_index)
}

@[keep_args_alive]
fn C.vkCreateIndirectCommandsLayoutNV(device Device, p_create_info &IndirectCommandsLayoutCreateInfoNV, p_allocator &AllocationCallbacks, p_indirect_commands_layout &IndirectCommandsLayoutNV) Result

pub type PFN_vkCreateIndirectCommandsLayoutNV = fn (device Device, p_create_info &IndirectCommandsLayoutCreateInfoNV, p_allocator &AllocationCallbacks, p_indirect_commands_layout &IndirectCommandsLayoutNV) Result

@[inline]
pub fn create_indirect_commands_layout_nv(device Device,
	p_create_info &IndirectCommandsLayoutCreateInfoNV,
	p_allocator &AllocationCallbacks,
	p_indirect_commands_layout &IndirectCommandsLayoutNV) Result {
	return C.vkCreateIndirectCommandsLayoutNV(device, p_create_info, p_allocator, p_indirect_commands_layout)
}

@[keep_args_alive]
fn C.vkDestroyIndirectCommandsLayoutNV(device Device, indirect_commands_layout IndirectCommandsLayoutNV, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyIndirectCommandsLayoutNV = fn (device Device, indirect_commands_layout IndirectCommandsLayoutNV, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_indirect_commands_layout_nv(device Device,
	indirect_commands_layout IndirectCommandsLayoutNV,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyIndirectCommandsLayoutNV(device, indirect_commands_layout, p_allocator)
}

pub const nv_inherited_viewport_scissor_spec_version = 1
pub const nv_inherited_viewport_scissor_extension_name = c'VK_NV_inherited_viewport_scissor'
// PhysicalDeviceInheritedViewportScissorFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceInheritedViewportScissorFeaturesNV = C.VkPhysicalDeviceInheritedViewportScissorFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceInheritedViewportScissorFeaturesNV {
pub mut:
	sType                      StructureType = StructureType.physical_device_inherited_viewport_scissor_features_nv
	pNext                      voidptr       = unsafe { nil }
	inheritedViewportScissor2D Bool32
}

// CommandBufferInheritanceViewportScissorInfoNV extends VkCommandBufferInheritanceInfo
pub type CommandBufferInheritanceViewportScissorInfoNV = C.VkCommandBufferInheritanceViewportScissorInfoNV

@[typedef]
pub struct C.VkCommandBufferInheritanceViewportScissorInfoNV {
pub mut:
	sType              StructureType = StructureType.command_buffer_inheritance_viewport_scissor_info_nv
	pNext              voidptr       = unsafe { nil }
	viewportScissor2D  Bool32
	viewportDepthCount u32
	pViewportDepths    &Viewport
}

pub const ext_texel_buffer_alignment_spec_version = 1
pub const ext_texel_buffer_alignment_extension_name = c'VK_EXT_texel_buffer_alignment'
// PhysicalDeviceTexelBufferAlignmentFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceTexelBufferAlignmentFeaturesEXT = C.VkPhysicalDeviceTexelBufferAlignmentFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceTexelBufferAlignmentFeaturesEXT {
pub mut:
	sType                StructureType = StructureType.physical_device_texel_buffer_alignment_features_ext
	pNext                voidptr       = unsafe { nil }
	texelBufferAlignment Bool32
}

pub type PhysicalDeviceTexelBufferAlignmentPropertiesEXT = C.VkPhysicalDeviceTexelBufferAlignmentProperties

pub const qcom_render_pass_transform_spec_version = 5
pub const qcom_render_pass_transform_extension_name = c'VK_QCOM_render_pass_transform'
// RenderPassTransformBeginInfoQCOM extends VkRenderPassBeginInfo
pub type RenderPassTransformBeginInfoQCOM = C.VkRenderPassTransformBeginInfoQCOM

@[typedef]
pub struct C.VkRenderPassTransformBeginInfoQCOM {
pub mut:
	sType     StructureType = StructureType.render_pass_transform_begin_info_qcom
	pNext     voidptr       = unsafe { nil }
	transform SurfaceTransformFlagBitsKHR
}

// CommandBufferInheritanceRenderPassTransformInfoQCOM extends VkCommandBufferInheritanceInfo
pub type CommandBufferInheritanceRenderPassTransformInfoQCOM = C.VkCommandBufferInheritanceRenderPassTransformInfoQCOM

@[typedef]
pub struct C.VkCommandBufferInheritanceRenderPassTransformInfoQCOM {
pub mut:
	sType      StructureType = StructureType.command_buffer_inheritance_render_pass_transform_info_qcom
	pNext      voidptr       = unsafe { nil }
	transform  SurfaceTransformFlagBitsKHR
	renderArea Rect2D
}

pub const ext_depth_bias_control_spec_version = 1
pub const ext_depth_bias_control_extension_name = c'VK_EXT_depth_bias_control'

pub enum DepthBiasRepresentationEXT as u32 {
	least_representable_value_format      = 0
	least_representable_value_force_unorm = 1
	float                                 = 2
	max_enum_ext                          = max_int
}
// PhysicalDeviceDepthBiasControlFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDepthBiasControlFeaturesEXT = C.VkPhysicalDeviceDepthBiasControlFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDepthBiasControlFeaturesEXT {
pub mut:
	sType                                           StructureType = StructureType.physical_device_depth_bias_control_features_ext
	pNext                                           voidptr       = unsafe { nil }
	depthBiasControl                                Bool32
	leastRepresentableValueForceUnormRepresentation Bool32
	floatRepresentation                             Bool32
	depthBiasExact                                  Bool32
}

pub type DepthBiasInfoEXT = C.VkDepthBiasInfoEXT

@[typedef]
pub struct C.VkDepthBiasInfoEXT {
pub mut:
	sType                   StructureType = StructureType.depth_bias_info_ext
	pNext                   voidptr       = unsafe { nil }
	depthBiasConstantFactor f32
	depthBiasClamp          f32
	depthBiasSlopeFactor    f32
}

// DepthBiasRepresentationInfoEXT extends VkDepthBiasInfoEXT,VkPipelineRasterizationStateCreateInfo
pub type DepthBiasRepresentationInfoEXT = C.VkDepthBiasRepresentationInfoEXT

@[typedef]
pub struct C.VkDepthBiasRepresentationInfoEXT {
pub mut:
	sType                   StructureType = StructureType.depth_bias_representation_info_ext
	pNext                   voidptr       = unsafe { nil }
	depthBiasRepresentation DepthBiasRepresentationEXT
	depthBiasExact          Bool32
}

@[keep_args_alive]
fn C.vkCmdSetDepthBias2EXT(command_buffer CommandBuffer, p_depth_bias_info &DepthBiasInfoEXT)

pub type PFN_vkCmdSetDepthBias2EXT = fn (command_buffer CommandBuffer, p_depth_bias_info &DepthBiasInfoEXT)

@[inline]
pub fn cmd_set_depth_bias2_ext(command_buffer CommandBuffer,
	p_depth_bias_info &DepthBiasInfoEXT) {
	C.vkCmdSetDepthBias2EXT(command_buffer, p_depth_bias_info)
}

pub const ext_device_memory_report_spec_version = 2
pub const ext_device_memory_report_extension_name = c'VK_EXT_device_memory_report'

pub enum DeviceMemoryReportEventTypeEXT as u32 {
	allocate          = 0
	free              = 1
	import            = 2
	unimport          = 3
	allocation_failed = 4
	max_enum_ext      = max_int
}
pub type DeviceMemoryReportFlagsEXT = u32

// PhysicalDeviceDeviceMemoryReportFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDeviceMemoryReportFeaturesEXT = C.VkPhysicalDeviceDeviceMemoryReportFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDeviceMemoryReportFeaturesEXT {
pub mut:
	sType              StructureType = StructureType.physical_device_device_memory_report_features_ext
	pNext              voidptr       = unsafe { nil }
	deviceMemoryReport Bool32
}

pub type DeviceMemoryReportCallbackDataEXT = C.VkDeviceMemoryReportCallbackDataEXT

@[typedef]
pub struct C.VkDeviceMemoryReportCallbackDataEXT {
pub mut:
	sType          StructureType = StructureType.device_memory_report_callback_data_ext
	pNext          voidptr       = unsafe { nil }
	flags          DeviceMemoryReportFlagsEXT
	type           DeviceMemoryReportEventTypeEXT
	memoryObjectId u64
	size           DeviceSize
	objectType     ObjectType
	objectHandle   u64
	heapIndex      u32
}

pub type PFN_vkDeviceMemoryReportCallbackEXT = fn (&DeviceMemoryReportCallbackDataEXT, voidptr)

// DeviceDeviceMemoryReportCreateInfoEXT extends VkDeviceCreateInfo
pub type DeviceDeviceMemoryReportCreateInfoEXT = C.VkDeviceDeviceMemoryReportCreateInfoEXT

@[typedef]
pub struct C.VkDeviceDeviceMemoryReportCreateInfoEXT {
pub mut:
	sType           StructureType = StructureType.device_device_memory_report_create_info_ext
	pNext           voidptr       = unsafe { nil }
	flags           DeviceMemoryReportFlagsEXT
	pfnUserCallback PFN_vkDeviceMemoryReportCallbackEXT = unsafe { nil }
	pUserData       voidptr = unsafe { nil }
}

pub const ext_acquire_drm_display_spec_version = 1
pub const ext_acquire_drm_display_extension_name = c'VK_EXT_acquire_drm_display'

@[keep_args_alive]
fn C.vkAcquireDrmDisplayEXT(physical_device PhysicalDevice, drm_fd i32, display DisplayKHR) Result

pub type PFN_vkAcquireDrmDisplayEXT = fn (physical_device PhysicalDevice, drm_fd i32, display DisplayKHR) Result

@[inline]
pub fn acquire_drm_display_ext(physical_device PhysicalDevice,
	drm_fd i32,
	display DisplayKHR) Result {
	return C.vkAcquireDrmDisplayEXT(physical_device, drm_fd, display)
}

@[keep_args_alive]
fn C.vkGetDrmDisplayEXT(physical_device PhysicalDevice, drm_fd i32, connector_id u32, display &DisplayKHR) Result

pub type PFN_vkGetDrmDisplayEXT = fn (physical_device PhysicalDevice, drm_fd i32, connector_id u32, display &DisplayKHR) Result

@[inline]
pub fn get_drm_display_ext(physical_device PhysicalDevice,
	drm_fd i32,
	connector_id u32,
	display &DisplayKHR) Result {
	return C.vkGetDrmDisplayEXT(physical_device, drm_fd, connector_id, display)
}

pub const ext_robustness_2_spec_version = 1
pub const ext_robustness_2_extension_name = c'VK_EXT_robustness2'

pub type PhysicalDeviceRobustness2FeaturesEXT = C.VkPhysicalDeviceRobustness2FeaturesKHR

pub type PhysicalDeviceRobustness2PropertiesEXT = C.VkPhysicalDeviceRobustness2PropertiesKHR

pub const ext_custom_border_color_spec_version = 12
pub const ext_custom_border_color_extension_name = c'VK_EXT_custom_border_color'
// SamplerCustomBorderColorCreateInfoEXT extends VkSamplerCreateInfo
pub type SamplerCustomBorderColorCreateInfoEXT = C.VkSamplerCustomBorderColorCreateInfoEXT

@[typedef]
pub struct C.VkSamplerCustomBorderColorCreateInfoEXT {
pub mut:
	sType             StructureType = StructureType.sampler_custom_border_color_create_info_ext
	pNext             voidptr       = unsafe { nil }
	customBorderColor ClearColorValue
	format            Format
}

// PhysicalDeviceCustomBorderColorPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceCustomBorderColorPropertiesEXT = C.VkPhysicalDeviceCustomBorderColorPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceCustomBorderColorPropertiesEXT {
pub mut:
	sType                        StructureType = StructureType.physical_device_custom_border_color_properties_ext
	pNext                        voidptr       = unsafe { nil }
	maxCustomBorderColorSamplers u32
}

// PhysicalDeviceCustomBorderColorFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCustomBorderColorFeaturesEXT = C.VkPhysicalDeviceCustomBorderColorFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceCustomBorderColorFeaturesEXT {
pub mut:
	sType                          StructureType = StructureType.physical_device_custom_border_color_features_ext
	pNext                          voidptr       = unsafe { nil }
	customBorderColors             Bool32
	customBorderColorWithoutFormat Bool32
}

pub const google_user_type_spec_version = 1
pub const google_user_type_extension_name = c'VK_GOOGE_user_type'

pub const nv_present_barrier_spec_version = 1
pub const nv_present_barrier_extension_name = c'VK_NV_present_barrier'
// PhysicalDevicePresentBarrierFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePresentBarrierFeaturesNV = C.VkPhysicalDevicePresentBarrierFeaturesNV

@[typedef]
pub struct C.VkPhysicalDevicePresentBarrierFeaturesNV {
pub mut:
	sType          StructureType = StructureType.physical_device_present_barrier_features_nv
	pNext          voidptr       = unsafe { nil }
	presentBarrier Bool32
}

// SurfaceCapabilitiesPresentBarrierNV extends VkSurfaceCapabilities2KHR
pub type SurfaceCapabilitiesPresentBarrierNV = C.VkSurfaceCapabilitiesPresentBarrierNV

@[typedef]
pub struct C.VkSurfaceCapabilitiesPresentBarrierNV {
pub mut:
	sType                   StructureType = StructureType.surface_capabilities_present_barrier_nv
	pNext                   voidptr       = unsafe { nil }
	presentBarrierSupported Bool32
}

// SwapchainPresentBarrierCreateInfoNV extends VkSwapchainCreateInfoKHR
pub type SwapchainPresentBarrierCreateInfoNV = C.VkSwapchainPresentBarrierCreateInfoNV

@[typedef]
pub struct C.VkSwapchainPresentBarrierCreateInfoNV {
pub mut:
	sType                StructureType = StructureType.swapchain_present_barrier_create_info_nv
	pNext                voidptr       = unsafe { nil }
	presentBarrierEnable Bool32
}

pub type PrivateDataSlotEXT = voidptr

pub const ext_private_data_spec_version = 1
pub const ext_private_data_extension_name = c'VK_EXT_private_data'

pub type PrivateDataSlotCreateFlagsEXT = u32
pub type PhysicalDevicePrivateDataFeaturesEXT = C.VkPhysicalDevicePrivateDataFeatures

pub type DevicePrivateDataCreateInfoEXT = C.VkDevicePrivateDataCreateInfo

pub type PrivateDataSlotCreateInfoEXT = C.VkPrivateDataSlotCreateInfo

@[keep_args_alive]
fn C.vkCreatePrivateDataSlotEXT(device Device, p_create_info &PrivateDataSlotCreateInfo, p_allocator &AllocationCallbacks, p_private_data_slot &PrivateDataSlot) Result

pub type PFN_vkCreatePrivateDataSlotEXT = fn (device Device, p_create_info &PrivateDataSlotCreateInfo, p_allocator &AllocationCallbacks, p_private_data_slot &PrivateDataSlot) Result

@[inline]
pub fn create_private_data_slot_ext(device Device,
	p_create_info &PrivateDataSlotCreateInfo,
	p_allocator &AllocationCallbacks,
	p_private_data_slot &PrivateDataSlot) Result {
	return C.vkCreatePrivateDataSlotEXT(device, p_create_info, p_allocator, p_private_data_slot)
}

@[keep_args_alive]
fn C.vkDestroyPrivateDataSlotEXT(device Device, private_data_slot PrivateDataSlot, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyPrivateDataSlotEXT = fn (device Device, private_data_slot PrivateDataSlot, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_private_data_slot_ext(device Device,
	private_data_slot PrivateDataSlot,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyPrivateDataSlotEXT(device, private_data_slot, p_allocator)
}

@[keep_args_alive]
fn C.vkSetPrivateDataEXT(device Device, object_type ObjectType, object_handle u64, private_data_slot PrivateDataSlot, data u64) Result

pub type PFN_vkSetPrivateDataEXT = fn (device Device, object_type ObjectType, object_handle u64, private_data_slot PrivateDataSlot, data u64) Result

@[inline]
pub fn set_private_data_ext(device Device,
	object_type ObjectType,
	object_handle u64,
	private_data_slot PrivateDataSlot,
	data u64) Result {
	return C.vkSetPrivateDataEXT(device, object_type, object_handle, private_data_slot,
		data)
}

@[keep_args_alive]
fn C.vkGetPrivateDataEXT(device Device, object_type ObjectType, object_handle u64, private_data_slot PrivateDataSlot, p_data &u64)

pub type PFN_vkGetPrivateDataEXT = fn (device Device, object_type ObjectType, object_handle u64, private_data_slot PrivateDataSlot, p_data &u64)

@[inline]
pub fn get_private_data_ext(device Device,
	object_type ObjectType,
	object_handle u64,
	private_data_slot PrivateDataSlot,
	p_data &u64) {
	C.vkGetPrivateDataEXT(device, object_type, object_handle, private_data_slot, p_data)
}

pub const ext_pipeline_creation_cache_control_spec_version = 3
pub const ext_pipeline_creation_cache_control_extension_name = c'VK_EXT_pipeline_creation_cache_control'

pub type PhysicalDevicePipelineCreationCacheControlFeaturesEXT = C.VkPhysicalDevicePipelineCreationCacheControlFeatures

pub const nv_device_diagnostics_config_spec_version = 2
pub const nv_device_diagnostics_config_extension_name = c'VK_NV_device_diagnostics_config'

pub enum DeviceDiagnosticsConfigFlagBitsNV as u32 {
	enable_shader_debug_info      = u32(0x00000001)
	enable_resource_tracking      = u32(0x00000002)
	enable_automatic_checkpoints  = u32(0x00000004)
	enable_shader_error_reporting = u32(0x00000008)
	max_enum_nv                   = max_int
}
pub type DeviceDiagnosticsConfigFlagsNV = u32

// PhysicalDeviceDiagnosticsConfigFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDiagnosticsConfigFeaturesNV = C.VkPhysicalDeviceDiagnosticsConfigFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceDiagnosticsConfigFeaturesNV {
pub mut:
	sType             StructureType = StructureType.physical_device_diagnostics_config_features_nv
	pNext             voidptr       = unsafe { nil }
	diagnosticsConfig Bool32
}

// DeviceDiagnosticsConfigCreateInfoNV extends VkDeviceCreateInfo
pub type DeviceDiagnosticsConfigCreateInfoNV = C.VkDeviceDiagnosticsConfigCreateInfoNV

@[typedef]
pub struct C.VkDeviceDiagnosticsConfigCreateInfoNV {
pub mut:
	sType StructureType = StructureType.device_diagnostics_config_create_info_nv
	pNext voidptr       = unsafe { nil }
	flags DeviceDiagnosticsConfigFlagsNV
}

pub const qcom_render_pass_store_ops_spec_version = 2
pub const qcom_render_pass_store_ops_extension_name = c'VK_QCOM_render_pass_store_ops'

// Pointer to VkCudaModuleNV_T
pub type CudaModuleNV = voidptr

// Pointer to VkCudaFunctionNV_T
pub type CudaFunctionNV = voidptr

pub const nv_cuda_kernel_launch_spec_version = 2
pub const nv_cuda_kernel_launch_extension_name = c'VK_NV_cuda_kernel_launch'

pub type CudaModuleCreateInfoNV = C.VkCudaModuleCreateInfoNV

@[typedef]
pub struct C.VkCudaModuleCreateInfoNV {
pub mut:
	sType    StructureType
	pNext    voidptr = unsafe { nil }
	dataSize usize
	pData    voidptr
}

pub type CudaFunctionCreateInfoNV = C.VkCudaFunctionCreateInfoNV

@[typedef]
pub struct C.VkCudaFunctionCreateInfoNV {
pub mut:
	sType  StructureType
	pNext  voidptr = unsafe { nil }
	module CudaModuleNV
	pName  &char
}

pub type CudaLaunchInfoNV = C.VkCudaLaunchInfoNV

@[typedef]
pub struct C.VkCudaLaunchInfoNV {
pub mut:
	sType          StructureType
	pNext          voidptr = unsafe { nil }
	function       CudaFunctionNV
	gridDimX       u32
	gridDimY       u32
	gridDimZ       u32
	blockDimX      u32
	blockDimY      u32
	blockDimZ      u32
	sharedMemBytes u32
	paramCount     usize
	pParams        &voidptr
	extraCount     usize
	pExtras        &voidptr
}

// PhysicalDeviceCudaKernelLaunchFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCudaKernelLaunchFeaturesNV = C.VkPhysicalDeviceCudaKernelLaunchFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceCudaKernelLaunchFeaturesNV {
pub mut:
	sType                    StructureType
	pNext                    voidptr = unsafe { nil }
	cudaKernelLaunchFeatures Bool32
}

// PhysicalDeviceCudaKernelLaunchPropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceCudaKernelLaunchPropertiesNV = C.VkPhysicalDeviceCudaKernelLaunchPropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceCudaKernelLaunchPropertiesNV {
pub mut:
	sType                  StructureType
	pNext                  voidptr = unsafe { nil }
	computeCapabilityMinor u32
	computeCapabilityMajor u32
}

@[keep_args_alive]
fn C.vkCreateCudaModuleNV(device Device, p_create_info &CudaModuleCreateInfoNV, p_allocator &AllocationCallbacks, p_module &CudaModuleNV) Result

pub type PFN_vkCreateCudaModuleNV = fn (device Device, p_create_info &CudaModuleCreateInfoNV, p_allocator &AllocationCallbacks, p_module &CudaModuleNV) Result

@[inline]
pub fn create_cuda_module_nv(device Device,
	p_create_info &CudaModuleCreateInfoNV,
	p_allocator &AllocationCallbacks,
	p_module &CudaModuleNV) Result {
	return C.vkCreateCudaModuleNV(device, p_create_info, p_allocator, p_module)
}

@[keep_args_alive]
fn C.vkGetCudaModuleCacheNV(device Device, vkmodule CudaModuleNV, p_cache_size &usize, p_cache_data voidptr) Result

pub type PFN_vkGetCudaModuleCacheNV = fn (device Device, vkmodule CudaModuleNV, p_cache_size &usize, p_cache_data voidptr) Result

@[inline]
pub fn get_cuda_module_cache_nv(device Device,
	vkmodule CudaModuleNV,
	p_cache_size &usize,
	p_cache_data voidptr) Result {
	return C.vkGetCudaModuleCacheNV(device, vkmodule, p_cache_size, p_cache_data)
}

@[keep_args_alive]
fn C.vkCreateCudaFunctionNV(device Device, p_create_info &CudaFunctionCreateInfoNV, p_allocator &AllocationCallbacks, p_function &CudaFunctionNV) Result

pub type PFN_vkCreateCudaFunctionNV = fn (device Device, p_create_info &CudaFunctionCreateInfoNV, p_allocator &AllocationCallbacks, p_function &CudaFunctionNV) Result

@[inline]
pub fn create_cuda_function_nv(device Device,
	p_create_info &CudaFunctionCreateInfoNV,
	p_allocator &AllocationCallbacks,
	p_function &CudaFunctionNV) Result {
	return C.vkCreateCudaFunctionNV(device, p_create_info, p_allocator, p_function)
}

@[keep_args_alive]
fn C.vkDestroyCudaModuleNV(device Device, vkmodule CudaModuleNV, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyCudaModuleNV = fn (device Device, vkmodule CudaModuleNV, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_cuda_module_nv(device Device,
	vkmodule CudaModuleNV,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyCudaModuleNV(device, vkmodule, p_allocator)
}

@[keep_args_alive]
fn C.vkDestroyCudaFunctionNV(device Device, function CudaFunctionNV, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyCudaFunctionNV = fn (device Device, function CudaFunctionNV, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_cuda_function_nv(device Device,
	function CudaFunctionNV,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyCudaFunctionNV(device, function, p_allocator)
}

@[keep_args_alive]
fn C.vkCmdCudaLaunchKernelNV(command_buffer CommandBuffer, p_launch_info &CudaLaunchInfoNV)

pub type PFN_vkCmdCudaLaunchKernelNV = fn (command_buffer CommandBuffer, p_launch_info &CudaLaunchInfoNV)

@[inline]
pub fn cmd_cuda_launch_kernel_nv(command_buffer CommandBuffer,
	p_launch_info &CudaLaunchInfoNV) {
	C.vkCmdCudaLaunchKernelNV(command_buffer, p_launch_info)
}

pub const qcom_tile_shading_spec_version = 2
pub const qcom_tile_shading_extension_name = c'VK_QCOM_tile_shading'

pub enum TileShadingRenderPassFlagBitsQCOM as u32 {
	enable             = u32(0x00000001)
	per_tile_execution = u32(0x00000002)
	max_enum_qcom      = max_int
}
pub type TileShadingRenderPassFlagsQCOM = u32

// PhysicalDeviceTileShadingFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceTileShadingFeaturesQCOM = C.VkPhysicalDeviceTileShadingFeaturesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceTileShadingFeaturesQCOM {
pub mut:
	sType                         StructureType = StructureType.physical_device_tile_shading_features_qcom
	pNext                         voidptr       = unsafe { nil }
	tileShading                   Bool32
	tileShadingFragmentStage      Bool32
	tileShadingColorAttachments   Bool32
	tileShadingDepthAttachments   Bool32
	tileShadingStencilAttachments Bool32
	tileShadingInputAttachments   Bool32
	tileShadingSampledAttachments Bool32
	tileShadingPerTileDraw        Bool32
	tileShadingPerTileDispatch    Bool32
	tileShadingDispatchTile       Bool32
	tileShadingApron              Bool32
	tileShadingAnisotropicApron   Bool32
	tileShadingAtomicOps          Bool32
	tileShadingImageProcessing    Bool32
}

// PhysicalDeviceTileShadingPropertiesQCOM extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceTileShadingPropertiesQCOM = C.VkPhysicalDeviceTileShadingPropertiesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceTileShadingPropertiesQCOM {
pub mut:
	sType              StructureType = StructureType.physical_device_tile_shading_properties_qcom
	pNext              voidptr       = unsafe { nil }
	maxApronSize       u32
	preferNonCoherent  Bool32
	tileGranularity    Extent2D
	maxTileShadingRate Extent2D
}

// RenderPassTileShadingCreateInfoQCOM extends VkRenderPassCreateInfo,VkRenderPassCreateInfo2,VkRenderingInfo,VkCommandBufferInheritanceInfo
pub type RenderPassTileShadingCreateInfoQCOM = C.VkRenderPassTileShadingCreateInfoQCOM

@[typedef]
pub struct C.VkRenderPassTileShadingCreateInfoQCOM {
pub mut:
	sType         StructureType = StructureType.render_pass_tile_shading_create_info_qcom
	pNext         voidptr       = unsafe { nil }
	flags         TileShadingRenderPassFlagsQCOM
	tileApronSize Extent2D
}

pub type PerTileBeginInfoQCOM = C.VkPerTileBeginInfoQCOM

@[typedef]
pub struct C.VkPerTileBeginInfoQCOM {
pub mut:
	sType StructureType = StructureType.per_tile_begin_info_qcom
	pNext voidptr       = unsafe { nil }
}

pub type PerTileEndInfoQCOM = C.VkPerTileEndInfoQCOM

@[typedef]
pub struct C.VkPerTileEndInfoQCOM {
pub mut:
	sType StructureType = StructureType.per_tile_end_info_qcom
	pNext voidptr       = unsafe { nil }
}

pub type DispatchTileInfoQCOM = C.VkDispatchTileInfoQCOM

@[typedef]
pub struct C.VkDispatchTileInfoQCOM {
pub mut:
	sType StructureType = StructureType.dispatch_tile_info_qcom
	pNext voidptr       = unsafe { nil }
}

@[keep_args_alive]
fn C.vkCmdDispatchTileQCOM(command_buffer CommandBuffer, p_dispatch_tile_info &DispatchTileInfoQCOM)

pub type PFN_vkCmdDispatchTileQCOM = fn (command_buffer CommandBuffer, p_dispatch_tile_info &DispatchTileInfoQCOM)

@[inline]
pub fn cmd_dispatch_tile_qcom(command_buffer CommandBuffer,
	p_dispatch_tile_info &DispatchTileInfoQCOM) {
	C.vkCmdDispatchTileQCOM(command_buffer, p_dispatch_tile_info)
}

@[keep_args_alive]
fn C.vkCmdBeginPerTileExecutionQCOM(command_buffer CommandBuffer, p_per_tile_begin_info &PerTileBeginInfoQCOM)

pub type PFN_vkCmdBeginPerTileExecutionQCOM = fn (command_buffer CommandBuffer, p_per_tile_begin_info &PerTileBeginInfoQCOM)

@[inline]
pub fn cmd_begin_per_tile_execution_qcom(command_buffer CommandBuffer,
	p_per_tile_begin_info &PerTileBeginInfoQCOM) {
	C.vkCmdBeginPerTileExecutionQCOM(command_buffer, p_per_tile_begin_info)
}

@[keep_args_alive]
fn C.vkCmdEndPerTileExecutionQCOM(command_buffer CommandBuffer, p_per_tile_end_info &PerTileEndInfoQCOM)

pub type PFN_vkCmdEndPerTileExecutionQCOM = fn (command_buffer CommandBuffer, p_per_tile_end_info &PerTileEndInfoQCOM)

@[inline]
pub fn cmd_end_per_tile_execution_qcom(command_buffer CommandBuffer,
	p_per_tile_end_info &PerTileEndInfoQCOM) {
	C.vkCmdEndPerTileExecutionQCOM(command_buffer, p_per_tile_end_info)
}

pub const nv_low_latency_spec_version = 1
pub const nv_low_latency_extension_name = c'VK_NV_low_latency'
// QueryLowLatencySupportNV extends VkSemaphoreCreateInfo
pub type QueryLowLatencySupportNV = C.VkQueryLowLatencySupportNV

@[typedef]
pub struct C.VkQueryLowLatencySupportNV {
pub mut:
	sType                  StructureType = StructureType.query_low_latency_support_nv
	pNext                  voidptr       = unsafe { nil }
	pQueriedLowLatencyData voidptr
}

// Pointer to VkAccelerationStructureKHR_T
pub type AccelerationStructureKHR = voidptr

pub const ext_descriptor_buffer_spec_version = 1
pub const ext_descriptor_buffer_extension_name = c'VK_EXT_descriptor_buffer'
// PhysicalDeviceDescriptorBufferPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceDescriptorBufferPropertiesEXT = C.VkPhysicalDeviceDescriptorBufferPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDescriptorBufferPropertiesEXT {
pub mut:
	sType                                                StructureType = StructureType.physical_device_descriptor_buffer_properties_ext
	pNext                                                voidptr       = unsafe { nil }
	combinedImageSamplerDescriptorSingleArray            Bool32
	bufferlessPushDescriptors                            Bool32
	allowSamplerImageViewPostSubmitCreation              Bool32
	descriptorBufferOffsetAlignment                      DeviceSize
	maxDescriptorBufferBindings                          u32
	maxResourceDescriptorBufferBindings                  u32
	maxSamplerDescriptorBufferBindings                   u32
	maxEmbeddedImmutableSamplerBindings                  u32
	maxEmbeddedImmutableSamplers                         u32
	bufferCaptureReplayDescriptorDataSize                usize
	imageCaptureReplayDescriptorDataSize                 usize
	imageViewCaptureReplayDescriptorDataSize             usize
	samplerCaptureReplayDescriptorDataSize               usize
	accelerationStructureCaptureReplayDescriptorDataSize usize
	samplerDescriptorSize                                usize
	combinedImageSamplerDescriptorSize                   usize
	sampledImageDescriptorSize                           usize
	storageImageDescriptorSize                           usize
	uniformTexelBufferDescriptorSize                     usize
	robustUniformTexelBufferDescriptorSize               usize
	storageTexelBufferDescriptorSize                     usize
	robustStorageTexelBufferDescriptorSize               usize
	uniformBufferDescriptorSize                          usize
	robustUniformBufferDescriptorSize                    usize
	storageBufferDescriptorSize                          usize
	robustStorageBufferDescriptorSize                    usize
	inputAttachmentDescriptorSize                        usize
	accelerationStructureDescriptorSize                  usize
	maxSamplerDescriptorBufferRange                      DeviceSize
	maxResourceDescriptorBufferRange                     DeviceSize
	samplerDescriptorBufferAddressSpaceSize              DeviceSize
	resourceDescriptorBufferAddressSpaceSize             DeviceSize
	descriptorBufferAddressSpaceSize                     DeviceSize
}

// PhysicalDeviceDescriptorBufferDensityMapPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceDescriptorBufferDensityMapPropertiesEXT = C.VkPhysicalDeviceDescriptorBufferDensityMapPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDescriptorBufferDensityMapPropertiesEXT {
pub mut:
	sType                                        StructureType = StructureType.physical_device_descriptor_buffer_density_map_properties_ext
	pNext                                        voidptr       = unsafe { nil }
	combinedImageSamplerDensityMapDescriptorSize usize
}

// PhysicalDeviceDescriptorBufferFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDescriptorBufferFeaturesEXT = C.VkPhysicalDeviceDescriptorBufferFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDescriptorBufferFeaturesEXT {
pub mut:
	sType                              StructureType = StructureType.physical_device_descriptor_buffer_features_ext
	pNext                              voidptr       = unsafe { nil }
	descriptorBuffer                   Bool32
	descriptorBufferCaptureReplay      Bool32
	descriptorBufferImageLayoutIgnored Bool32
	descriptorBufferPushDescriptors    Bool32
}

pub type DescriptorAddressInfoEXT = C.VkDescriptorAddressInfoEXT

@[typedef]
pub struct C.VkDescriptorAddressInfoEXT {
pub mut:
	sType   StructureType = StructureType.descriptor_address_info_ext
	pNext   voidptr       = unsafe { nil }
	address DeviceAddress
	range   DeviceSize
	format  Format
}

pub type DescriptorBufferBindingInfoEXT = C.VkDescriptorBufferBindingInfoEXT

@[typedef]
pub struct C.VkDescriptorBufferBindingInfoEXT {
pub mut:
	sType   StructureType = StructureType.descriptor_buffer_binding_info_ext
	pNext   voidptr       = unsafe { nil }
	address DeviceAddress
	usage   BufferUsageFlags
}

// DescriptorBufferBindingPushDescriptorBufferHandleEXT extends VkDescriptorBufferBindingInfoEXT
pub type DescriptorBufferBindingPushDescriptorBufferHandleEXT = C.VkDescriptorBufferBindingPushDescriptorBufferHandleEXT

@[typedef]
pub struct C.VkDescriptorBufferBindingPushDescriptorBufferHandleEXT {
pub mut:
	sType  StructureType = StructureType.descriptor_buffer_binding_push_descriptor_buffer_handle_ext
	pNext  voidptr       = unsafe { nil }
	buffer Buffer
}

pub type DescriptorDataEXT = C.VkDescriptorDataEXT

@[typedef]
pub union C.VkDescriptorDataEXT {
pub mut:
	pSampler              &Sampler
	pCombinedImageSampler &DescriptorImageInfo
	pInputAttachmentImage &DescriptorImageInfo
	pSampledImage         &DescriptorImageInfo
	pStorageImage         &DescriptorImageInfo
	pUniformTexelBuffer   &DescriptorAddressInfoEXT
	pStorageTexelBuffer   &DescriptorAddressInfoEXT
	pUniformBuffer        &DescriptorAddressInfoEXT
	pStorageBuffer        &DescriptorAddressInfoEXT
	accelerationStructure DeviceAddress
}

pub type DescriptorGetInfoEXT = C.VkDescriptorGetInfoEXT

@[typedef]
pub struct C.VkDescriptorGetInfoEXT {
pub mut:
	sType StructureType = StructureType.descriptor_get_info_ext
	pNext voidptr       = unsafe { nil }
	type  DescriptorType
	data  DescriptorDataEXT
}

pub type BufferCaptureDescriptorDataInfoEXT = C.VkBufferCaptureDescriptorDataInfoEXT

@[typedef]
pub struct C.VkBufferCaptureDescriptorDataInfoEXT {
pub mut:
	sType  StructureType = StructureType.buffer_capture_descriptor_data_info_ext
	pNext  voidptr       = unsafe { nil }
	buffer Buffer
}

pub type ImageCaptureDescriptorDataInfoEXT = C.VkImageCaptureDescriptorDataInfoEXT

@[typedef]
pub struct C.VkImageCaptureDescriptorDataInfoEXT {
pub mut:
	sType StructureType = StructureType.image_capture_descriptor_data_info_ext
	pNext voidptr       = unsafe { nil }
	image Image
}

pub type ImageViewCaptureDescriptorDataInfoEXT = C.VkImageViewCaptureDescriptorDataInfoEXT

@[typedef]
pub struct C.VkImageViewCaptureDescriptorDataInfoEXT {
pub mut:
	sType     StructureType = StructureType.image_view_capture_descriptor_data_info_ext
	pNext     voidptr       = unsafe { nil }
	imageView ImageView
}

pub type SamplerCaptureDescriptorDataInfoEXT = C.VkSamplerCaptureDescriptorDataInfoEXT

@[typedef]
pub struct C.VkSamplerCaptureDescriptorDataInfoEXT {
pub mut:
	sType   StructureType = StructureType.sampler_capture_descriptor_data_info_ext
	pNext   voidptr       = unsafe { nil }
	sampler Sampler
}

// OpaqueCaptureDescriptorDataCreateInfoEXT extends VkBufferCreateInfo,VkImageCreateInfo,VkImageViewCreateInfo,VkSamplerCreateInfo,VkAccelerationStructureCreateInfoKHR,VkAccelerationStructureCreateInfoNV,VkTensorCreateInfoARM,VkTensorViewCreateInfoARM
pub type OpaqueCaptureDescriptorDataCreateInfoEXT = C.VkOpaqueCaptureDescriptorDataCreateInfoEXT

@[typedef]
pub struct C.VkOpaqueCaptureDescriptorDataCreateInfoEXT {
pub mut:
	sType                       StructureType = StructureType.opaque_capture_descriptor_data_create_info_ext
	pNext                       voidptr       = unsafe { nil }
	opaqueCaptureDescriptorData voidptr
}

pub type AccelerationStructureCaptureDescriptorDataInfoEXT = C.VkAccelerationStructureCaptureDescriptorDataInfoEXT

@[typedef]
pub struct C.VkAccelerationStructureCaptureDescriptorDataInfoEXT {
pub mut:
	sType                   StructureType = StructureType.acceleration_structure_capture_descriptor_data_info_ext
	pNext                   voidptr       = unsafe { nil }
	accelerationStructure   AccelerationStructureKHR
	accelerationStructureNV AccelerationStructureNV
}

@[keep_args_alive]
fn C.vkGetDescriptorSetLayoutSizeEXT(device Device, layout DescriptorSetLayout, p_layout_size_in_bytes &DeviceSize)

pub type PFN_vkGetDescriptorSetLayoutSizeEXT = fn (device Device, layout DescriptorSetLayout, p_layout_size_in_bytes &DeviceSize)

@[inline]
pub fn get_descriptor_set_layout_size_ext(device Device,
	layout DescriptorSetLayout,
	p_layout_size_in_bytes &DeviceSize) {
	C.vkGetDescriptorSetLayoutSizeEXT(device, layout, p_layout_size_in_bytes)
}

@[keep_args_alive]
fn C.vkGetDescriptorSetLayoutBindingOffsetEXT(device Device, layout DescriptorSetLayout, binding u32, p_offset &DeviceSize)

pub type PFN_vkGetDescriptorSetLayoutBindingOffsetEXT = fn (device Device, layout DescriptorSetLayout, binding u32, p_offset &DeviceSize)

@[inline]
pub fn get_descriptor_set_layout_binding_offset_ext(device Device,
	layout DescriptorSetLayout,
	binding u32,
	p_offset &DeviceSize) {
	C.vkGetDescriptorSetLayoutBindingOffsetEXT(device, layout, binding, p_offset)
}

@[keep_args_alive]
fn C.vkGetDescriptorEXT(device Device, p_descriptor_info &DescriptorGetInfoEXT, data_size usize, p_descriptor voidptr)

pub type PFN_vkGetDescriptorEXT = fn (device Device, p_descriptor_info &DescriptorGetInfoEXT, data_size usize, p_descriptor voidptr)

@[inline]
pub fn get_descriptor_ext(device Device,
	p_descriptor_info &DescriptorGetInfoEXT,
	data_size usize,
	p_descriptor voidptr) {
	C.vkGetDescriptorEXT(device, p_descriptor_info, data_size, p_descriptor)
}

@[keep_args_alive]
fn C.vkCmdBindDescriptorBuffersEXT(command_buffer CommandBuffer, buffer_count u32, p_binding_infos &DescriptorBufferBindingInfoEXT)

pub type PFN_vkCmdBindDescriptorBuffersEXT = fn (command_buffer CommandBuffer, buffer_count u32, p_binding_infos &DescriptorBufferBindingInfoEXT)

@[inline]
pub fn cmd_bind_descriptor_buffers_ext(command_buffer CommandBuffer,
	buffer_count u32,
	p_binding_infos &DescriptorBufferBindingInfoEXT) {
	C.vkCmdBindDescriptorBuffersEXT(command_buffer, buffer_count, p_binding_infos)
}

@[keep_args_alive]
fn C.vkCmdSetDescriptorBufferOffsetsEXT(command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, layout PipelineLayout, first_set u32, set_count u32, p_buffer_indices &u32, p_offsets &DeviceSize)

pub type PFN_vkCmdSetDescriptorBufferOffsetsEXT = fn (command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, layout PipelineLayout, first_set u32, set_count u32, p_buffer_indices &u32, p_offsets &DeviceSize)

@[inline]
pub fn cmd_set_descriptor_buffer_offsets_ext(command_buffer CommandBuffer,
	pipeline_bind_point PipelineBindPoint,
	layout PipelineLayout,
	first_set u32,
	set_count u32,
	p_buffer_indices &u32,
	p_offsets &DeviceSize) {
	C.vkCmdSetDescriptorBufferOffsetsEXT(command_buffer, pipeline_bind_point, layout,
		first_set, set_count, p_buffer_indices, p_offsets)
}

@[keep_args_alive]
fn C.vkCmdBindDescriptorBufferEmbeddedSamplersEXT(command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, layout PipelineLayout, set u32)

pub type PFN_vkCmdBindDescriptorBufferEmbeddedSamplersEXT = fn (command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, layout PipelineLayout, set u32)

@[inline]
pub fn cmd_bind_descriptor_buffer_embedded_samplers_ext(command_buffer CommandBuffer,
	pipeline_bind_point PipelineBindPoint,
	layout PipelineLayout,
	set u32) {
	C.vkCmdBindDescriptorBufferEmbeddedSamplersEXT(command_buffer, pipeline_bind_point,
		layout, set)
}

@[keep_args_alive]
fn C.vkGetBufferOpaqueCaptureDescriptorDataEXT(device Device, p_info &BufferCaptureDescriptorDataInfoEXT, p_data voidptr) Result

pub type PFN_vkGetBufferOpaqueCaptureDescriptorDataEXT = fn (device Device, p_info &BufferCaptureDescriptorDataInfoEXT, p_data voidptr) Result

@[inline]
pub fn get_buffer_opaque_capture_descriptor_data_ext(device Device,
	p_info &BufferCaptureDescriptorDataInfoEXT,
	p_data voidptr) Result {
	return C.vkGetBufferOpaqueCaptureDescriptorDataEXT(device, p_info, p_data)
}

@[keep_args_alive]
fn C.vkGetImageOpaqueCaptureDescriptorDataEXT(device Device, p_info &ImageCaptureDescriptorDataInfoEXT, p_data voidptr) Result

pub type PFN_vkGetImageOpaqueCaptureDescriptorDataEXT = fn (device Device, p_info &ImageCaptureDescriptorDataInfoEXT, p_data voidptr) Result

@[inline]
pub fn get_image_opaque_capture_descriptor_data_ext(device Device,
	p_info &ImageCaptureDescriptorDataInfoEXT,
	p_data voidptr) Result {
	return C.vkGetImageOpaqueCaptureDescriptorDataEXT(device, p_info, p_data)
}

@[keep_args_alive]
fn C.vkGetImageViewOpaqueCaptureDescriptorDataEXT(device Device, p_info &ImageViewCaptureDescriptorDataInfoEXT, p_data voidptr) Result

pub type PFN_vkGetImageViewOpaqueCaptureDescriptorDataEXT = fn (device Device, p_info &ImageViewCaptureDescriptorDataInfoEXT, p_data voidptr) Result

@[inline]
pub fn get_image_view_opaque_capture_descriptor_data_ext(device Device,
	p_info &ImageViewCaptureDescriptorDataInfoEXT,
	p_data voidptr) Result {
	return C.vkGetImageViewOpaqueCaptureDescriptorDataEXT(device, p_info, p_data)
}

@[keep_args_alive]
fn C.vkGetSamplerOpaqueCaptureDescriptorDataEXT(device Device, p_info &SamplerCaptureDescriptorDataInfoEXT, p_data voidptr) Result

pub type PFN_vkGetSamplerOpaqueCaptureDescriptorDataEXT = fn (device Device, p_info &SamplerCaptureDescriptorDataInfoEXT, p_data voidptr) Result

@[inline]
pub fn get_sampler_opaque_capture_descriptor_data_ext(device Device,
	p_info &SamplerCaptureDescriptorDataInfoEXT,
	p_data voidptr) Result {
	return C.vkGetSamplerOpaqueCaptureDescriptorDataEXT(device, p_info, p_data)
}

@[keep_args_alive]
fn C.vkGetAccelerationStructureOpaqueCaptureDescriptorDataEXT(device Device, p_info &AccelerationStructureCaptureDescriptorDataInfoEXT, p_data voidptr) Result

pub type PFN_vkGetAccelerationStructureOpaqueCaptureDescriptorDataEXT = fn (device Device, p_info &AccelerationStructureCaptureDescriptorDataInfoEXT, p_data voidptr) Result

@[inline]
pub fn get_acceleration_structure_opaque_capture_descriptor_data_ext(device Device,
	p_info &AccelerationStructureCaptureDescriptorDataInfoEXT,
	p_data voidptr) Result {
	return C.vkGetAccelerationStructureOpaqueCaptureDescriptorDataEXT(device, p_info,
		p_data)
}

pub const ext_graphics_pipeline_library_spec_version = 1
pub const ext_graphics_pipeline_library_extension_name = c'VK_EXT_graphics_pipeline_library'

pub enum GraphicsPipelineLibraryFlagBitsEXT as u32 {
	vertex_input_interface    = u32(0x00000001)
	pre_rasterization_shaders = u32(0x00000002)
	fragment_shader           = u32(0x00000004)
	fragment_output_interface = u32(0x00000008)
	max_enum_ext              = max_int
}
pub type GraphicsPipelineLibraryFlagsEXT = u32

// PhysicalDeviceGraphicsPipelineLibraryFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceGraphicsPipelineLibraryFeaturesEXT = C.VkPhysicalDeviceGraphicsPipelineLibraryFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceGraphicsPipelineLibraryFeaturesEXT {
pub mut:
	sType                   StructureType = StructureType.physical_device_graphics_pipeline_library_features_ext
	pNext                   voidptr       = unsafe { nil }
	graphicsPipelineLibrary Bool32
}

// PhysicalDeviceGraphicsPipelineLibraryPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceGraphicsPipelineLibraryPropertiesEXT = C.VkPhysicalDeviceGraphicsPipelineLibraryPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceGraphicsPipelineLibraryPropertiesEXT {
pub mut:
	sType                                                     StructureType = StructureType.physical_device_graphics_pipeline_library_properties_ext
	pNext                                                     voidptr       = unsafe { nil }
	graphicsPipelineLibraryFastLinking                        Bool32
	graphicsPipelineLibraryIndependentInterpolationDecoration Bool32
}

// GraphicsPipelineLibraryCreateInfoEXT extends VkGraphicsPipelineCreateInfo
pub type GraphicsPipelineLibraryCreateInfoEXT = C.VkGraphicsPipelineLibraryCreateInfoEXT

@[typedef]
pub struct C.VkGraphicsPipelineLibraryCreateInfoEXT {
pub mut:
	sType StructureType = StructureType.graphics_pipeline_library_create_info_ext
	pNext voidptr       = unsafe { nil }
	flags GraphicsPipelineLibraryFlagsEXT
}

pub const amd_shader_early_and_late_fragment_tests_spec_version = 1
pub const amd_shader_early_and_late_fragment_tests_extension_name = c'VK_AMD_shader_early_and_late_fragment_tests'
// PhysicalDeviceShaderEarlyAndLateFragmentTestsFeaturesAMD extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderEarlyAndLateFragmentTestsFeaturesAMD = C.VkPhysicalDeviceShaderEarlyAndLateFragmentTestsFeaturesAMD

@[typedef]
pub struct C.VkPhysicalDeviceShaderEarlyAndLateFragmentTestsFeaturesAMD {
pub mut:
	sType                           StructureType = StructureType.physical_device_shader_early_and_late_fragment_tests_features_amd
	pNext                           voidptr       = unsafe { nil }
	shaderEarlyAndLateFragmentTests Bool32
}

pub const nv_fragment_shading_rate_enums_spec_version = 1
pub const nv_fragment_shading_rate_enums_extension_name = c'VK_NV_fragment_shading_rate_enums'

pub enum FragmentShadingRateTypeNV as u32 {
	fragment_size = 0
	enums         = 1
	max_enum_nv   = max_int
}

pub enum FragmentShadingRateNV as u32 {
	_1_invocation_per_pixel     = 0
	_1_invocation_per1x2_pixels = 1
	_1_invocation_per2x1_pixels = 4
	_1_invocation_per2x2_pixels = 5
	_1_invocation_per2x4_pixels = 6
	_1_invocation_per4x2_pixels = 9
	_1_invocation_per4x4_pixels = 10
	_2_invocations_per_pixel    = 11
	_4_invocations_per_pixel    = 12
	_8_invocations_per_pixel    = 13
	_16_invocations_per_pixel   = 14
	no_invocations              = 15
	max_enum_nv                 = max_int
}
// PhysicalDeviceFragmentShadingRateEnumsFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceFragmentShadingRateEnumsFeaturesNV = C.VkPhysicalDeviceFragmentShadingRateEnumsFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceFragmentShadingRateEnumsFeaturesNV {
pub mut:
	sType                            StructureType = StructureType.physical_device_fragment_shading_rate_enums_features_nv
	pNext                            voidptr       = unsafe { nil }
	fragmentShadingRateEnums         Bool32
	supersampleFragmentShadingRates  Bool32
	noInvocationFragmentShadingRates Bool32
}

// PhysicalDeviceFragmentShadingRateEnumsPropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceFragmentShadingRateEnumsPropertiesNV = C.VkPhysicalDeviceFragmentShadingRateEnumsPropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceFragmentShadingRateEnumsPropertiesNV {
pub mut:
	sType                                 StructureType = StructureType.physical_device_fragment_shading_rate_enums_properties_nv
	pNext                                 voidptr       = unsafe { nil }
	maxFragmentShadingRateInvocationCount SampleCountFlagBits
}

// PipelineFragmentShadingRateEnumStateCreateInfoNV extends VkGraphicsPipelineCreateInfo
pub type PipelineFragmentShadingRateEnumStateCreateInfoNV = C.VkPipelineFragmentShadingRateEnumStateCreateInfoNV

@[typedef]
pub struct C.VkPipelineFragmentShadingRateEnumStateCreateInfoNV {
pub mut:
	sType           StructureType = StructureType.pipeline_fragment_shading_rate_enum_state_create_info_nv
	pNext           voidptr       = unsafe { nil }
	shadingRateType FragmentShadingRateTypeNV
	shadingRate     FragmentShadingRateNV
	combinerOps     [2]FragmentShadingRateCombinerOpKHR
}

/*@[keep_args_alive]
fn C.vkCmdSetFragmentShadingRateEnumNV(
 command_buffer CommandBuffer,  shading_rate FragmentShadingRateNV,  combiner_ops [2]FragmentShadingRateCombinerOpKHR)
pub type PFN_vkCmdSetFragmentShadingRateEnumNV = fn(command_buffer CommandBuffer, shading_rate FragmentShadingRateNV, combiner_ops [2]FragmentShadingRateCombinerOpKHR)
@[inline]
pub fn cmd_set_fragment_shading_rate_enum_nv(
command_buffer CommandBuffer,
shading_rate FragmentShadingRateNV,
combiner_ops [2]FragmentShadingRateCombinerOpKHR) {
    C.vkCmdSetFragmentShadingRateEnumNV( command_buffer, shading_rate, combiner_ops)
}

*/

pub const nv_ray_tracing_motion_blur_spec_version = 1
pub const nv_ray_tracing_motion_blur_extension_name = c'VK_NV_ray_tracing_motion_blur'

pub enum AccelerationStructureMotionInstanceTypeNV as u32 {
	static        = 0
	matrix_motion = 1
	srt_motion    = 2
	max_enum_nv   = max_int
}
pub type AccelerationStructureMotionInfoFlagsNV = u32
pub type AccelerationStructureMotionInstanceFlagsNV = u32
pub type DeviceOrHostAddressConstKHR = C.VkDeviceOrHostAddressConstKHR

@[typedef]
pub union C.VkDeviceOrHostAddressConstKHR {
pub mut:
	deviceAddress DeviceAddress
	hostAddress   voidptr
}

// AccelerationStructureGeometryMotionTrianglesDataNV extends VkAccelerationStructureGeometryTrianglesDataKHR
pub type AccelerationStructureGeometryMotionTrianglesDataNV = C.VkAccelerationStructureGeometryMotionTrianglesDataNV

@[typedef]
pub struct C.VkAccelerationStructureGeometryMotionTrianglesDataNV {
pub mut:
	sType      StructureType = StructureType.acceleration_structure_geometry_motion_triangles_data_nv
	pNext      voidptr       = unsafe { nil }
	vertexData DeviceOrHostAddressConstKHR
}

// AccelerationStructureMotionInfoNV extends VkAccelerationStructureCreateInfoKHR
pub type AccelerationStructureMotionInfoNV = C.VkAccelerationStructureMotionInfoNV

@[typedef]
pub struct C.VkAccelerationStructureMotionInfoNV {
pub mut:
	sType        StructureType = StructureType.acceleration_structure_motion_info_nv
	pNext        voidptr       = unsafe { nil }
	maxInstances u32
	flags        AccelerationStructureMotionInfoFlagsNV
}

pub type AccelerationStructureMatrixMotionInstanceNV = C.VkAccelerationStructureMatrixMotionInstanceNV

@[typedef]
pub struct C.VkAccelerationStructureMatrixMotionInstanceNV {
pub mut:
	transformT0                            TransformMatrixKHR
	transformT1                            TransformMatrixKHR
	instanceCustomIndex                    u32
	mask                                   u32
	instanceShaderBindingTableRecordOffset u32
	flags                                  GeometryInstanceFlagsKHR
	accelerationStructureReference         u64
}

pub type SRTDataNV = C.VkSRTDataNV

@[typedef]
pub struct C.VkSRTDataNV {
pub mut:
	sx  f32
	a   f32
	b   f32
	pvx f32
	sy  f32
	c   f32
	pvy f32
	sz  f32
	pvz f32
	qx  f32
	qy  f32
	qz  f32
	qw  f32
	tx  f32
	ty  f32
	tz  f32
}

pub type AccelerationStructureSRTMotionInstanceNV = C.VkAccelerationStructureSRTMotionInstanceNV

@[typedef]
pub struct C.VkAccelerationStructureSRTMotionInstanceNV {
pub mut:
	transformT0                            SRTDataNV
	transformT1                            SRTDataNV
	instanceCustomIndex                    u32
	mask                                   u32
	instanceShaderBindingTableRecordOffset u32
	flags                                  GeometryInstanceFlagsKHR
	accelerationStructureReference         u64
}

pub type AccelerationStructureMotionInstanceDataNV = C.VkAccelerationStructureMotionInstanceDataNV

@[typedef]
pub union C.VkAccelerationStructureMotionInstanceDataNV {
pub mut:
	staticInstance       AccelerationStructureInstanceKHR
	matrixMotionInstance AccelerationStructureMatrixMotionInstanceNV
	srtMotionInstance    AccelerationStructureSRTMotionInstanceNV
}

pub type AccelerationStructureMotionInstanceNV = C.VkAccelerationStructureMotionInstanceNV

@[typedef]
pub struct C.VkAccelerationStructureMotionInstanceNV {
pub mut:
	type  AccelerationStructureMotionInstanceTypeNV
	flags AccelerationStructureMotionInstanceFlagsNV
	data  AccelerationStructureMotionInstanceDataNV
}

// PhysicalDeviceRayTracingMotionBlurFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRayTracingMotionBlurFeaturesNV = C.VkPhysicalDeviceRayTracingMotionBlurFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceRayTracingMotionBlurFeaturesNV {
pub mut:
	sType                                         StructureType = StructureType.physical_device_ray_tracing_motion_blur_features_nv
	pNext                                         voidptr       = unsafe { nil }
	rayTracingMotionBlur                          Bool32
	rayTracingMotionBlurPipelineTraceRaysIndirect Bool32
}

pub const ext_ycbcr_2plane_444_formats_spec_version = 1
pub const ext_ycbcr_2plane_444_formats_extension_name = c'VK_EXT_ycbcr_2plane_444_formats'
// PhysicalDeviceYcbcr2Plane444FormatsFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceYcbcr2Plane444FormatsFeaturesEXT = C.VkPhysicalDeviceYcbcr2Plane444FormatsFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceYcbcr2Plane444FormatsFeaturesEXT {
pub mut:
	sType                 StructureType = StructureType.physical_device_ycbcr2_plane444_formats_features_ext
	pNext                 voidptr       = unsafe { nil }
	ycbcr2plane444Formats Bool32
}

pub const ext_fragment_density_map_2_spec_version = 1
pub const ext_fragment_density_map_2_extension_name = c'VK_EXT_fragment_density_map2'
// PhysicalDeviceFragmentDensityMap2FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceFragmentDensityMap2FeaturesEXT = C.VkPhysicalDeviceFragmentDensityMap2FeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceFragmentDensityMap2FeaturesEXT {
pub mut:
	sType                      StructureType = StructureType.physical_device_fragment_density_map2_features_ext
	pNext                      voidptr       = unsafe { nil }
	fragmentDensityMapDeferred Bool32
}

// PhysicalDeviceFragmentDensityMap2PropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceFragmentDensityMap2PropertiesEXT = C.VkPhysicalDeviceFragmentDensityMap2PropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceFragmentDensityMap2PropertiesEXT {
pub mut:
	sType                                     StructureType = StructureType.physical_device_fragment_density_map2_properties_ext
	pNext                                     voidptr       = unsafe { nil }
	subsampledLoads                           Bool32
	subsampledCoarseReconstructionEarlyAccess Bool32
	maxSubsampledArrayLayers                  u32
	maxDescriptorSetSubsampledSamplers        u32
}

pub const qcom_rotated_copy_commands_spec_version = 2
pub const qcom_rotated_copy_commands_extension_name = c'VK_QCOM_rotated_copy_commands'
// CopyCommandTransformInfoQCOM extends VkBufferImageCopy2,VkImageBlit2
pub type CopyCommandTransformInfoQCOM = C.VkCopyCommandTransformInfoQCOM

@[typedef]
pub struct C.VkCopyCommandTransformInfoQCOM {
pub mut:
	sType     StructureType = StructureType.copy_command_transform_info_qcom
	pNext     voidptr       = unsafe { nil }
	transform SurfaceTransformFlagBitsKHR
}

pub const ext_image_robustness_spec_version = 1
pub const ext_image_robustness_extension_name = c'VK_EXT_image_robustness'

pub type PhysicalDeviceImageRobustnessFeaturesEXT = C.VkPhysicalDeviceImageRobustnessFeatures

pub const ext_image_compression_control_spec_version = 1
pub const ext_image_compression_control_extension_name = c'VK_EXT_image_compression_control'

pub enum ImageCompressionFlagBitsEXT as u32 {
	default             = 0
	fixed_rate_default  = u32(0x00000001)
	fixed_rate_explicit = u32(0x00000002)
	disabled            = u32(0x00000004)
	max_enum_ext        = max_int
}
pub type ImageCompressionFlagsEXT = u32

pub enum ImageCompressionFixedRateFlagBitsEXT as u32 {
	none         = 0
	_1bpc        = u32(0x00000001)
	_2bpc        = u32(0x00000002)
	_3bpc        = u32(0x00000004)
	_4bpc        = u32(0x00000008)
	_5bpc        = u32(0x00000010)
	_6bpc        = u32(0x00000020)
	_7bpc        = u32(0x00000040)
	_8bpc        = u32(0x00000080)
	_9bpc        = u32(0x00000100)
	_10bpc       = u32(0x00000200)
	_11bpc       = u32(0x00000400)
	_12bpc       = u32(0x00000800)
	_13bpc       = u32(0x00001000)
	_14bpc       = u32(0x00002000)
	_15bpc       = u32(0x00004000)
	_16bpc       = u32(0x00008000)
	_17bpc       = u32(0x00010000)
	_18bpc       = u32(0x00020000)
	_19bpc       = u32(0x00040000)
	_20bpc       = u32(0x00080000)
	_21bpc       = u32(0x00100000)
	_22bpc       = u32(0x00200000)
	_23bpc       = u32(0x00400000)
	_24bpc       = u32(0x00800000)
	max_enum_ext = max_int
}
pub type ImageCompressionFixedRateFlagsEXT = u32

// PhysicalDeviceImageCompressionControlFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceImageCompressionControlFeaturesEXT = C.VkPhysicalDeviceImageCompressionControlFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceImageCompressionControlFeaturesEXT {
pub mut:
	sType                   StructureType = StructureType.physical_device_image_compression_control_features_ext
	pNext                   voidptr       = unsafe { nil }
	imageCompressionControl Bool32
}

// ImageCompressionControlEXT extends VkImageCreateInfo,VkSwapchainCreateInfoKHR,VkPhysicalDeviceImageFormatInfo2
pub type ImageCompressionControlEXT = C.VkImageCompressionControlEXT

@[typedef]
pub struct C.VkImageCompressionControlEXT {
pub mut:
	sType                        StructureType = StructureType.image_compression_control_ext
	pNext                        voidptr       = unsafe { nil }
	flags                        ImageCompressionFlagsEXT
	compressionControlPlaneCount u32
	pFixedRateFlags              &ImageCompressionFixedRateFlagsEXT
}

// ImageCompressionPropertiesEXT extends VkImageFormatProperties2,VkSurfaceFormat2KHR,VkSubresourceLayout2
pub type ImageCompressionPropertiesEXT = C.VkImageCompressionPropertiesEXT

@[typedef]
pub struct C.VkImageCompressionPropertiesEXT {
pub mut:
	sType                          StructureType = StructureType.image_compression_properties_ext
	pNext                          voidptr       = unsafe { nil }
	imageCompressionFlags          ImageCompressionFlagsEXT
	imageCompressionFixedRateFlags ImageCompressionFixedRateFlagsEXT
}

pub const ext_attachment_feedback_loop_layout_spec_version = 2
pub const ext_attachment_feedback_loop_layout_extension_name = c'VK_EXT_attachment_feedback_loop_layout'
// PhysicalDeviceAttachmentFeedbackLoopLayoutFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceAttachmentFeedbackLoopLayoutFeaturesEXT = C.VkPhysicalDeviceAttachmentFeedbackLoopLayoutFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceAttachmentFeedbackLoopLayoutFeaturesEXT {
pub mut:
	sType                        StructureType = StructureType.physical_device_attachment_feedback_loop_layout_features_ext
	pNext                        voidptr       = unsafe { nil }
	attachmentFeedbackLoopLayout Bool32
}

pub const ext_4444_formats_spec_version = 1
pub const ext_4444_formats_extension_name = c'VK_EXT_4444_formats'
// PhysicalDevice4444FormatsFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevice4444FormatsFeaturesEXT = C.VkPhysicalDevice4444FormatsFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDevice4444FormatsFeaturesEXT {
pub mut:
	sType          StructureType = StructureType.physical_device4444_formats_features_ext
	pNext          voidptr       = unsafe { nil }
	formatA4R4G4B4 Bool32
	formatA4B4G4R4 Bool32
}

pub const ext_device_fault_spec_version = 2
pub const ext_device_fault_extension_name = c'VK_EXT_device_fault'

pub enum DeviceFaultAddressTypeEXT as u32 {
	none                        = 0
	read_invalid                = 1
	write_invalid               = 2
	execute_invalid             = 3
	instruction_pointer_unknown = 4
	instruction_pointer_invalid = 5
	instruction_pointer_fault   = 6
	max_enum_ext                = max_int
}

pub enum DeviceFaultVendorBinaryHeaderVersionEXT as u32 {
	one          = 1
	max_enum_ext = max_int
}
// PhysicalDeviceFaultFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceFaultFeaturesEXT = C.VkPhysicalDeviceFaultFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceFaultFeaturesEXT {
pub mut:
	sType                   StructureType = StructureType.physical_device_fault_features_ext
	pNext                   voidptr       = unsafe { nil }
	deviceFault             Bool32
	deviceFaultVendorBinary Bool32
}

pub type DeviceFaultCountsEXT = C.VkDeviceFaultCountsEXT

@[typedef]
pub struct C.VkDeviceFaultCountsEXT {
pub mut:
	sType            StructureType = StructureType.device_fault_counts_ext
	pNext            voidptr       = unsafe { nil }
	addressInfoCount u32
	vendorInfoCount  u32
	vendorBinarySize DeviceSize
}

pub type DeviceFaultAddressInfoEXT = C.VkDeviceFaultAddressInfoEXT

@[typedef]
pub struct C.VkDeviceFaultAddressInfoEXT {
pub mut:
	addressType      DeviceFaultAddressTypeEXT
	reportedAddress  DeviceAddress
	addressPrecision DeviceSize
}

pub type DeviceFaultVendorInfoEXT = C.VkDeviceFaultVendorInfoEXT

@[typedef]
pub struct C.VkDeviceFaultVendorInfoEXT {
pub mut:
	description     [max_description_size]char
	vendorFaultCode u64
	vendorFaultData u64
}

pub type DeviceFaultInfoEXT = C.VkDeviceFaultInfoEXT

@[typedef]
pub struct C.VkDeviceFaultInfoEXT {
pub mut:
	sType             StructureType = StructureType.device_fault_info_ext
	pNext             voidptr       = unsafe { nil }
	description       [max_description_size]char
	pAddressInfos     &DeviceFaultAddressInfoEXT
	pVendorInfos      &DeviceFaultVendorInfoEXT
	pVendorBinaryData voidptr
}

pub type DeviceFaultVendorBinaryHeaderVersionOneEXT = C.VkDeviceFaultVendorBinaryHeaderVersionOneEXT

@[typedef]
pub struct C.VkDeviceFaultVendorBinaryHeaderVersionOneEXT {
pub mut:
	headerSize            u32
	headerVersion         DeviceFaultVendorBinaryHeaderVersionEXT
	vendorID              u32
	deviceID              u32
	driverVersion         u32
	pipelineCacheUUID     [uuid_size]u8
	applicationNameOffset u32
	applicationVersion    u32
	engineNameOffset      u32
	engineVersion         u32
	apiVersion            u32
}

@[keep_args_alive]
fn C.vkGetDeviceFaultInfoEXT(device Device, mut p_fault_counts DeviceFaultCountsEXT, mut p_fault_info DeviceFaultInfoEXT) Result

pub type PFN_vkGetDeviceFaultInfoEXT = fn (device Device, mut p_fault_counts DeviceFaultCountsEXT, mut p_fault_info DeviceFaultInfoEXT) Result

@[inline]
pub fn get_device_fault_info_ext(device Device,
	mut p_fault_counts DeviceFaultCountsEXT,
	mut p_fault_info DeviceFaultInfoEXT) Result {
	return C.vkGetDeviceFaultInfoEXT(device, mut p_fault_counts, mut p_fault_info)
}

pub const arm_rasterization_order_attachment_access_spec_version = 1
pub const arm_rasterization_order_attachment_access_extension_name = c'VK_ARM_rasterization_order_attachment_access'
// PhysicalDeviceRasterizationOrderAttachmentAccessFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRasterizationOrderAttachmentAccessFeaturesEXT = C.VkPhysicalDeviceRasterizationOrderAttachmentAccessFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceRasterizationOrderAttachmentAccessFeaturesEXT {
pub mut:
	sType                                     StructureType = StructureType.physical_device_rasterization_order_attachment_access_features_ext
	pNext                                     voidptr       = unsafe { nil }
	rasterizationOrderColorAttachmentAccess   Bool32
	rasterizationOrderDepthAttachmentAccess   Bool32
	rasterizationOrderStencilAttachmentAccess Bool32
}

pub type PhysicalDeviceRasterizationOrderAttachmentAccessFeaturesARM = C.VkPhysicalDeviceRasterizationOrderAttachmentAccessFeaturesEXT

pub const ext_rgba10x6_formats_spec_version = 1
pub const ext_rgba10x6_formats_extension_name = c'VK_EXT_rgba10x6_formats'
// PhysicalDeviceRGBA10X6FormatsFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRGBA10X6FormatsFeaturesEXT = C.VkPhysicalDeviceRGBA10X6FormatsFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceRGBA10X6FormatsFeaturesEXT {
pub mut:
	sType                             StructureType = StructureType.physical_device_rgba10x6_formats_features_ext
	pNext                             voidptr       = unsafe { nil }
	formatRgba10x6WithoutYCbCrSampler Bool32
}

pub const valve_mutable_descriptor_type_spec_version = 1
pub const valve_mutable_descriptor_type_extension_name = c'VK_VAVE_mutable_descriptor_type'
// PhysicalDeviceMutableDescriptorTypeFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMutableDescriptorTypeFeaturesEXT = C.VkPhysicalDeviceMutableDescriptorTypeFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMutableDescriptorTypeFeaturesEXT {
pub mut:
	sType                 StructureType = StructureType.physical_device_mutable_descriptor_type_features_ext
	pNext                 voidptr       = unsafe { nil }
	mutableDescriptorType Bool32
}

pub type PhysicalDeviceMutableDescriptorTypeFeaturesVALVE = C.VkPhysicalDeviceMutableDescriptorTypeFeaturesEXT

pub type MutableDescriptorTypeListEXT = C.VkMutableDescriptorTypeListEXT

@[typedef]
pub struct C.VkMutableDescriptorTypeListEXT {
pub mut:
	descriptorTypeCount u32
	pDescriptorTypes    &DescriptorType
}

pub type MutableDescriptorTypeListVALVE = C.VkMutableDescriptorTypeListEXT

// MutableDescriptorTypeCreateInfoEXT extends VkDescriptorSetLayoutCreateInfo,VkDescriptorPoolCreateInfo
pub type MutableDescriptorTypeCreateInfoEXT = C.VkMutableDescriptorTypeCreateInfoEXT

@[typedef]
pub struct C.VkMutableDescriptorTypeCreateInfoEXT {
pub mut:
	sType                          StructureType = StructureType.mutable_descriptor_type_create_info_ext
	pNext                          voidptr       = unsafe { nil }
	mutableDescriptorTypeListCount u32
	pMutableDescriptorTypeLists    &MutableDescriptorTypeListEXT
}

pub type MutableDescriptorTypeCreateInfoVALVE = C.VkMutableDescriptorTypeCreateInfoEXT

pub const ext_vertex_input_dynamic_state_spec_version = 2
pub const ext_vertex_input_dynamic_state_extension_name = c'VK_EXT_vertex_input_dynamic_state'
// PhysicalDeviceVertexInputDynamicStateFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVertexInputDynamicStateFeaturesEXT = C.VkPhysicalDeviceVertexInputDynamicStateFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceVertexInputDynamicStateFeaturesEXT {
pub mut:
	sType                   StructureType = StructureType.physical_device_vertex_input_dynamic_state_features_ext
	pNext                   voidptr       = unsafe { nil }
	vertexInputDynamicState Bool32
}

pub type VertexInputBindingDescription2EXT = C.VkVertexInputBindingDescription2EXT

@[typedef]
pub struct C.VkVertexInputBindingDescription2EXT {
pub mut:
	sType     StructureType = StructureType.vertex_input_binding_description2_ext
	pNext     voidptr       = unsafe { nil }
	binding   u32
	stride    u32
	inputRate VertexInputRate
	divisor   u32
}

pub type VertexInputAttributeDescription2EXT = C.VkVertexInputAttributeDescription2EXT

@[typedef]
pub struct C.VkVertexInputAttributeDescription2EXT {
pub mut:
	sType    StructureType = StructureType.vertex_input_attribute_description2_ext
	pNext    voidptr       = unsafe { nil }
	location u32
	binding  u32
	format   Format
	offset   u32
}

@[keep_args_alive]
fn C.vkCmdSetVertexInputEXT(command_buffer CommandBuffer, vertex_binding_description_count u32, p_vertex_binding_descriptions &VertexInputBindingDescription2EXT, vertex_attribute_description_count u32, p_vertex_attribute_descriptions &VertexInputAttributeDescription2EXT)

pub type PFN_vkCmdSetVertexInputEXT = fn (command_buffer CommandBuffer, vertex_binding_description_count u32, p_vertex_binding_descriptions &VertexInputBindingDescription2EXT, vertex_attribute_description_count u32, p_vertex_attribute_descriptions &VertexInputAttributeDescription2EXT)

@[inline]
pub fn cmd_set_vertex_input_ext(command_buffer CommandBuffer,
	vertex_binding_description_count u32,
	p_vertex_binding_descriptions &VertexInputBindingDescription2EXT,
	vertex_attribute_description_count u32,
	p_vertex_attribute_descriptions &VertexInputAttributeDescription2EXT) {
	C.vkCmdSetVertexInputEXT(command_buffer, vertex_binding_description_count, p_vertex_binding_descriptions,
		vertex_attribute_description_count, p_vertex_attribute_descriptions)
}

pub const ext_physical_device_drm_spec_version = 1
pub const ext_physical_device_drm_extension_name = c'VK_EXT_physical_device_drm'
// PhysicalDeviceDrmPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceDrmPropertiesEXT = C.VkPhysicalDeviceDrmPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDrmPropertiesEXT {
pub mut:
	sType        StructureType = StructureType.physical_device_drm_properties_ext
	pNext        voidptr       = unsafe { nil }
	hasPrimary   Bool32
	hasRender    Bool32
	primaryMajor i64
	primaryMinor i64
	renderMajor  i64
	renderMinor  i64
}

pub const ext_device_address_binding_report_spec_version = 1
pub const ext_device_address_binding_report_extension_name = c'VK_EXT_device_address_binding_report'

pub enum DeviceAddressBindingTypeEXT as u32 {
	bind         = 0
	unbind       = 1
	max_enum_ext = max_int
}

pub enum DeviceAddressBindingFlagBitsEXT as u32 {
	internal_object = u32(0x00000001)
	max_enum_ext    = max_int
}
pub type DeviceAddressBindingFlagsEXT = u32

// PhysicalDeviceAddressBindingReportFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceAddressBindingReportFeaturesEXT = C.VkPhysicalDeviceAddressBindingReportFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceAddressBindingReportFeaturesEXT {
pub mut:
	sType                StructureType = StructureType.physical_device_address_binding_report_features_ext
	pNext                voidptr       = unsafe { nil }
	reportAddressBinding Bool32
}

// DeviceAddressBindingCallbackDataEXT extends VkDebugUtilsMessengerCallbackDataEXT
pub type DeviceAddressBindingCallbackDataEXT = C.VkDeviceAddressBindingCallbackDataEXT

@[typedef]
pub struct C.VkDeviceAddressBindingCallbackDataEXT {
pub mut:
	sType       StructureType = StructureType.device_address_binding_callback_data_ext
	pNext       voidptr       = unsafe { nil }
	flags       DeviceAddressBindingFlagsEXT
	baseAddress DeviceAddress
	size        DeviceSize
	bindingType DeviceAddressBindingTypeEXT
}

pub const ext_depth_clip_control_spec_version = 1
pub const ext_depth_clip_control_extension_name = c'VK_EXT_depth_clip_control'
// PhysicalDeviceDepthClipControlFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDepthClipControlFeaturesEXT = C.VkPhysicalDeviceDepthClipControlFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDepthClipControlFeaturesEXT {
pub mut:
	sType            StructureType = StructureType.physical_device_depth_clip_control_features_ext
	pNext            voidptr       = unsafe { nil }
	depthClipControl Bool32
}

// PipelineViewportDepthClipControlCreateInfoEXT extends VkPipelineViewportStateCreateInfo
pub type PipelineViewportDepthClipControlCreateInfoEXT = C.VkPipelineViewportDepthClipControlCreateInfoEXT

@[typedef]
pub struct C.VkPipelineViewportDepthClipControlCreateInfoEXT {
pub mut:
	sType            StructureType = StructureType.pipeline_viewport_depth_clip_control_create_info_ext
	pNext            voidptr       = unsafe { nil }
	negativeOneToOne Bool32
}

pub const ext_primitive_topology_list_restart_spec_version = 1
pub const ext_primitive_topology_list_restart_extension_name = c'VK_EXT_primitive_topology_list_restart'
// PhysicalDevicePrimitiveTopologyListRestartFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePrimitiveTopologyListRestartFeaturesEXT = C.VkPhysicalDevicePrimitiveTopologyListRestartFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDevicePrimitiveTopologyListRestartFeaturesEXT {
pub mut:
	sType                             StructureType = StructureType.physical_device_primitive_topology_list_restart_features_ext
	pNext                             voidptr       = unsafe { nil }
	primitiveTopologyListRestart      Bool32
	primitiveTopologyPatchListRestart Bool32
}

pub const ext_present_mode_fifo_latest_ready_spec_version = 1
pub const ext_present_mode_fifo_latest_ready_extension_name = c'VK_EXT_present_mode_fifo_latest_ready'

pub type PhysicalDevicePresentModeFifoLatestReadyFeaturesEXT = C.VkPhysicalDevicePresentModeFifoLatestReadyFeaturesKHR

pub const huawei_subpass_shading_spec_version = 3
pub const huawei_subpass_shading_extension_name = c'VK_HAWEI_subpass_shading'
// SubpassShadingPipelineCreateInfoHUAWEI extends VkComputePipelineCreateInfo
pub type SubpassShadingPipelineCreateInfoHUAWEI = C.VkSubpassShadingPipelineCreateInfoHUAWEI

@[typedef]
pub struct C.VkSubpassShadingPipelineCreateInfoHUAWEI {
pub mut:
	sType      StructureType = StructureType.subpass_shading_pipeline_create_info_huawei
	pNext      voidptr       = unsafe { nil }
	renderPass RenderPass
	subpass    u32
}

// PhysicalDeviceSubpassShadingFeaturesHUAWEI extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceSubpassShadingFeaturesHUAWEI = C.VkPhysicalDeviceSubpassShadingFeaturesHUAWEI

@[typedef]
pub struct C.VkPhysicalDeviceSubpassShadingFeaturesHUAWEI {
pub mut:
	sType          StructureType = StructureType.physical_device_subpass_shading_features_huawei
	pNext          voidptr       = unsafe { nil }
	subpassShading Bool32
}

// PhysicalDeviceSubpassShadingPropertiesHUAWEI extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceSubpassShadingPropertiesHUAWEI = C.VkPhysicalDeviceSubpassShadingPropertiesHUAWEI

@[typedef]
pub struct C.VkPhysicalDeviceSubpassShadingPropertiesHUAWEI {
pub mut:
	sType                                     StructureType = StructureType.physical_device_subpass_shading_properties_huawei
	pNext                                     voidptr       = unsafe { nil }
	maxSubpassShadingWorkgroupSizeAspectRatio u32
}

@[keep_args_alive]
fn C.vkGetDeviceSubpassShadingMaxWorkgroupSizeHUAWEI(device Device, renderpass RenderPass, mut p_max_workgroup_size Extent2D) Result

pub type PFN_vkGetDeviceSubpassShadingMaxWorkgroupSizeHUAWEI = fn (device Device, renderpass RenderPass, mut p_max_workgroup_size Extent2D) Result

@[inline]
pub fn get_device_subpass_shading_max_workgroup_size_huawei(device Device,
	renderpass RenderPass,
	mut p_max_workgroup_size Extent2D) Result {
	return C.vkGetDeviceSubpassShadingMaxWorkgroupSizeHUAWEI(device, renderpass, mut p_max_workgroup_size)
}

@[keep_args_alive]
fn C.vkCmdSubpassShadingHUAWEI(command_buffer CommandBuffer)

pub type PFN_vkCmdSubpassShadingHUAWEI = fn (command_buffer CommandBuffer)

@[inline]
pub fn cmd_subpass_shading_huawei(command_buffer CommandBuffer) {
	C.vkCmdSubpassShadingHUAWEI(command_buffer)
}

pub const huawei_invocation_mask_spec_version = 1
pub const huawei_invocation_mask_extension_name = c'VK_HAWEI_invocation_mask'
// PhysicalDeviceInvocationMaskFeaturesHUAWEI extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceInvocationMaskFeaturesHUAWEI = C.VkPhysicalDeviceInvocationMaskFeaturesHUAWEI

@[typedef]
pub struct C.VkPhysicalDeviceInvocationMaskFeaturesHUAWEI {
pub mut:
	sType          StructureType = StructureType.physical_device_invocation_mask_features_huawei
	pNext          voidptr       = unsafe { nil }
	invocationMask Bool32
}

@[keep_args_alive]
fn C.vkCmdBindInvocationMaskHUAWEI(command_buffer CommandBuffer, image_view ImageView, image_layout ImageLayout)

pub type PFN_vkCmdBindInvocationMaskHUAWEI = fn (command_buffer CommandBuffer, image_view ImageView, image_layout ImageLayout)

@[inline]
pub fn cmd_bind_invocation_mask_huawei(command_buffer CommandBuffer,
	image_view ImageView,
	image_layout ImageLayout) {
	C.vkCmdBindInvocationMaskHUAWEI(command_buffer, image_view, image_layout)
}

pub type RemoteAddressNV = voidptr

pub const nv_external_memory_rdma_spec_version = 1
pub const nv_external_memory_rdma_extension_name = c'VK_NV_external_memory_rdma'

pub type MemoryGetRemoteAddressInfoNV = C.VkMemoryGetRemoteAddressInfoNV

@[typedef]
pub struct C.VkMemoryGetRemoteAddressInfoNV {
pub mut:
	sType      StructureType = StructureType.memory_get_remote_address_info_nv
	pNext      voidptr       = unsafe { nil }
	memory     DeviceMemory
	handleType ExternalMemoryHandleTypeFlagBits
}

// PhysicalDeviceExternalMemoryRDMAFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceExternalMemoryRDMAFeaturesNV = C.VkPhysicalDeviceExternalMemoryRDMAFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceExternalMemoryRDMAFeaturesNV {
pub mut:
	sType              StructureType = StructureType.physical_device_external_memory_rdma_features_nv
	pNext              voidptr       = unsafe { nil }
	externalMemoryRDMA Bool32
}

@[keep_args_alive]
fn C.vkGetMemoryRemoteAddressNV(device Device, p_memory_get_remote_address_info &MemoryGetRemoteAddressInfoNV, p_address &RemoteAddressNV) Result

pub type PFN_vkGetMemoryRemoteAddressNV = fn (device Device, p_memory_get_remote_address_info &MemoryGetRemoteAddressInfoNV, p_address &RemoteAddressNV) Result

@[inline]
pub fn get_memory_remote_address_nv(device Device,
	p_memory_get_remote_address_info &MemoryGetRemoteAddressInfoNV,
	p_address &RemoteAddressNV) Result {
	return C.vkGetMemoryRemoteAddressNV(device, p_memory_get_remote_address_info, p_address)
}

pub const ext_pipeline_properties_spec_version = 1
pub const ext_pipeline_properties_extension_name = c'VK_EXT_pipeline_properties'

pub type PipelineInfoEXT = C.VkPipelineInfoKHR

pub type PipelinePropertiesIdentifierEXT = C.VkPipelinePropertiesIdentifierEXT

@[typedef]
pub struct C.VkPipelinePropertiesIdentifierEXT {
pub mut:
	sType              StructureType = StructureType.pipeline_properties_identifier_ext
	pNext              voidptr       = unsafe { nil }
	pipelineIdentifier [uuid_size]u8
}

// PhysicalDevicePipelinePropertiesFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePipelinePropertiesFeaturesEXT = C.VkPhysicalDevicePipelinePropertiesFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDevicePipelinePropertiesFeaturesEXT {
pub mut:
	sType                        StructureType = StructureType.physical_device_pipeline_properties_features_ext
	pNext                        voidptr       = unsafe { nil }
	pipelinePropertiesIdentifier Bool32
}

@[keep_args_alive]
fn C.vkGetPipelinePropertiesEXT(device Device, p_pipeline_info &PipelineInfoEXT, mut p_pipeline_properties BaseOutStructure) Result

pub type PFN_vkGetPipelinePropertiesEXT = fn (device Device, p_pipeline_info &PipelineInfoEXT, mut p_pipeline_properties BaseOutStructure) Result

@[inline]
pub fn get_pipeline_properties_ext(device Device,
	p_pipeline_info &PipelineInfoEXT,
	mut p_pipeline_properties BaseOutStructure) Result {
	return C.vkGetPipelinePropertiesEXT(device, p_pipeline_info, mut p_pipeline_properties)
}

pub const ext_frame_boundary_spec_version = 1
pub const ext_frame_boundary_extension_name = c'VK_EXT_frame_boundary'

pub enum FrameBoundaryFlagBitsEXT as u32 {
	frame_end    = u32(0x00000001)
	max_enum_ext = max_int
}
pub type FrameBoundaryFlagsEXT = u32

// PhysicalDeviceFrameBoundaryFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceFrameBoundaryFeaturesEXT = C.VkPhysicalDeviceFrameBoundaryFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceFrameBoundaryFeaturesEXT {
pub mut:
	sType         StructureType = StructureType.physical_device_frame_boundary_features_ext
	pNext         voidptr       = unsafe { nil }
	frameBoundary Bool32
}

// FrameBoundaryEXT extends VkSubmitInfo,VkSubmitInfo2,VkPresentInfoKHR,VkBindSparseInfo
pub type FrameBoundaryEXT = C.VkFrameBoundaryEXT

@[typedef]
pub struct C.VkFrameBoundaryEXT {
pub mut:
	sType       StructureType = StructureType.frame_boundary_ext
	pNext       voidptr       = unsafe { nil }
	flags       FrameBoundaryFlagsEXT
	frameID     u64
	imageCount  u32
	pImages     &Image
	bufferCount u32
	pBuffers    &Buffer
	tagName     u64
	tagSize     usize
	pTag        voidptr
}

pub const ext_multisampled_render_to_single_sampled_spec_version = 1
pub const ext_multisampled_render_to_single_sampled_extension_name = c'VK_EXT_multisampled_render_to_single_sampled'
// PhysicalDeviceMultisampledRenderToSingleSampledFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMultisampledRenderToSingleSampledFeaturesEXT = C.VkPhysicalDeviceMultisampledRenderToSingleSampledFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMultisampledRenderToSingleSampledFeaturesEXT {
pub mut:
	sType                             StructureType = StructureType.physical_device_multisampled_render_to_single_sampled_features_ext
	pNext                             voidptr       = unsafe { nil }
	multisampledRenderToSingleSampled Bool32
}

// SubpassResolvePerformanceQueryEXT extends VkFormatProperties2
pub type SubpassResolvePerformanceQueryEXT = C.VkSubpassResolvePerformanceQueryEXT

@[typedef]
pub struct C.VkSubpassResolvePerformanceQueryEXT {
pub mut:
	sType   StructureType = StructureType.subpass_resolve_performance_query_ext
	pNext   voidptr       = unsafe { nil }
	optimal Bool32
}

// MultisampledRenderToSingleSampledInfoEXT extends VkSubpassDescription2,VkRenderingInfo
pub type MultisampledRenderToSingleSampledInfoEXT = C.VkMultisampledRenderToSingleSampledInfoEXT

@[typedef]
pub struct C.VkMultisampledRenderToSingleSampledInfoEXT {
pub mut:
	sType                                   StructureType = StructureType.multisampled_render_to_single_sampled_info_ext
	pNext                                   voidptr       = unsafe { nil }
	multisampledRenderToSingleSampledEnable Bool32
	rasterizationSamples                    SampleCountFlagBits
}

pub const ext_extended_dynamic_state_2_spec_version = 1
pub const ext_extended_dynamic_state_2_extension_name = c'VK_EXT_extended_dynamic_state2'
// PhysicalDeviceExtendedDynamicState2FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceExtendedDynamicState2FeaturesEXT = C.VkPhysicalDeviceExtendedDynamicState2FeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceExtendedDynamicState2FeaturesEXT {
pub mut:
	sType                                   StructureType = StructureType.physical_device_extended_dynamic_state2_features_ext
	pNext                                   voidptr       = unsafe { nil }
	extendedDynamicState2                   Bool32
	extendedDynamicState2LogicOp            Bool32
	extendedDynamicState2PatchControlPoints Bool32
}

@[keep_args_alive]
fn C.vkCmdSetPatchControlPointsEXT(command_buffer CommandBuffer, patch_control_points u32)

pub type PFN_vkCmdSetPatchControlPointsEXT = fn (command_buffer CommandBuffer, patch_control_points u32)

@[inline]
pub fn cmd_set_patch_control_points_ext(command_buffer CommandBuffer,
	patch_control_points u32) {
	C.vkCmdSetPatchControlPointsEXT(command_buffer, patch_control_points)
}

@[keep_args_alive]
fn C.vkCmdSetRasterizerDiscardEnableEXT(command_buffer CommandBuffer, rasterizer_discard_enable Bool32)

pub type PFN_vkCmdSetRasterizerDiscardEnableEXT = fn (command_buffer CommandBuffer, rasterizer_discard_enable Bool32)

@[inline]
pub fn cmd_set_rasterizer_discard_enable_ext(command_buffer CommandBuffer,
	rasterizer_discard_enable Bool32) {
	C.vkCmdSetRasterizerDiscardEnableEXT(command_buffer, rasterizer_discard_enable)
}

@[keep_args_alive]
fn C.vkCmdSetDepthBiasEnableEXT(command_buffer CommandBuffer, depth_bias_enable Bool32)

pub type PFN_vkCmdSetDepthBiasEnableEXT = fn (command_buffer CommandBuffer, depth_bias_enable Bool32)

@[inline]
pub fn cmd_set_depth_bias_enable_ext(command_buffer CommandBuffer,
	depth_bias_enable Bool32) {
	C.vkCmdSetDepthBiasEnableEXT(command_buffer, depth_bias_enable)
}

@[keep_args_alive]
fn C.vkCmdSetLogicOpEXT(command_buffer CommandBuffer, logic_op LogicOp)

pub type PFN_vkCmdSetLogicOpEXT = fn (command_buffer CommandBuffer, logic_op LogicOp)

@[inline]
pub fn cmd_set_logic_op_ext(command_buffer CommandBuffer,
	logic_op LogicOp) {
	C.vkCmdSetLogicOpEXT(command_buffer, logic_op)
}

@[keep_args_alive]
fn C.vkCmdSetPrimitiveRestartEnableEXT(command_buffer CommandBuffer, primitive_restart_enable Bool32)

pub type PFN_vkCmdSetPrimitiveRestartEnableEXT = fn (command_buffer CommandBuffer, primitive_restart_enable Bool32)

@[inline]
pub fn cmd_set_primitive_restart_enable_ext(command_buffer CommandBuffer,
	primitive_restart_enable Bool32) {
	C.vkCmdSetPrimitiveRestartEnableEXT(command_buffer, primitive_restart_enable)
}

pub const ext_color_write_enable_spec_version = 1
pub const ext_color_write_enable_extension_name = c'VK_EXT_color_write_enable'
// PhysicalDeviceColorWriteEnableFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceColorWriteEnableFeaturesEXT = C.VkPhysicalDeviceColorWriteEnableFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceColorWriteEnableFeaturesEXT {
pub mut:
	sType            StructureType = StructureType.physical_device_color_write_enable_features_ext
	pNext            voidptr       = unsafe { nil }
	colorWriteEnable Bool32
}

// PipelineColorWriteCreateInfoEXT extends VkPipelineColorBlendStateCreateInfo
pub type PipelineColorWriteCreateInfoEXT = C.VkPipelineColorWriteCreateInfoEXT

@[typedef]
pub struct C.VkPipelineColorWriteCreateInfoEXT {
pub mut:
	sType              StructureType = StructureType.pipeline_color_write_create_info_ext
	pNext              voidptr       = unsafe { nil }
	attachmentCount    u32
	pColorWriteEnables &Bool32
}

@[keep_args_alive]
fn C.vkCmdSetColorWriteEnableEXT(command_buffer CommandBuffer, attachment_count u32, p_color_write_enables &Bool32)

pub type PFN_vkCmdSetColorWriteEnableEXT = fn (command_buffer CommandBuffer, attachment_count u32, p_color_write_enables &Bool32)

@[inline]
pub fn cmd_set_color_write_enable_ext(command_buffer CommandBuffer,
	attachment_count u32,
	p_color_write_enables &Bool32) {
	C.vkCmdSetColorWriteEnableEXT(command_buffer, attachment_count, p_color_write_enables)
}

pub const ext_primitives_generated_query_spec_version = 1
pub const ext_primitives_generated_query_extension_name = c'VK_EXT_primitives_generated_query'
// PhysicalDevicePrimitivesGeneratedQueryFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePrimitivesGeneratedQueryFeaturesEXT = C.VkPhysicalDevicePrimitivesGeneratedQueryFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDevicePrimitivesGeneratedQueryFeaturesEXT {
pub mut:
	sType                                         StructureType = StructureType.physical_device_primitives_generated_query_features_ext
	pNext                                         voidptr       = unsafe { nil }
	primitivesGeneratedQuery                      Bool32
	primitivesGeneratedQueryWithRasterizerDiscard Bool32
	primitivesGeneratedQueryWithNonZeroStreams    Bool32
}

pub const ext_global_priority_query_spec_version = 1
pub const ext_global_priority_query_extension_name = c'VK_EXT_global_priority_query'
pub const max_global_priority_size_ext = max_global_priority_size

pub type PhysicalDeviceGlobalPriorityQueryFeaturesEXT = C.VkPhysicalDeviceGlobalPriorityQueryFeatures

pub type QueueFamilyGlobalPriorityPropertiesEXT = C.VkQueueFamilyGlobalPriorityProperties

pub const valve_video_encode_rgb_conversion_spec_version = 1
pub const valve_video_encode_rgb_conversion_extension_name = c'VK_VAVE_video_encode_rgb_conversion'

pub enum VideoEncodeRgbModelConversionFlagBitsVALVE as u32 {
	rgb_identity   = u32(0x00000001)
	ycbcr_identity = u32(0x00000002)
	ycbcr709       = u32(0x00000004)
	ycbcr601       = u32(0x00000008)
	ycbcr2020      = u32(0x00000010)
	max_enum_valve = max_int
}
pub type VideoEncodeRgbModelConversionFlagsVALVE = u32

pub enum VideoEncodeRgbRangeCompressionFlagBitsVALVE as u32 {
	full_range     = u32(0x00000001)
	narrow_range   = u32(0x00000002)
	max_enum_valve = max_int
}
pub type VideoEncodeRgbRangeCompressionFlagsVALVE = u32

pub enum VideoEncodeRgbChromaOffsetFlagBitsVALVE as u32 {
	cosited_even   = u32(0x00000001)
	midpoint       = u32(0x00000002)
	max_enum_valve = max_int
}
pub type VideoEncodeRgbChromaOffsetFlagsVALVE = u32

// PhysicalDeviceVideoEncodeRgbConversionFeaturesVALVE extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVideoEncodeRgbConversionFeaturesVALVE = C.VkPhysicalDeviceVideoEncodeRgbConversionFeaturesVALVE

@[typedef]
pub struct C.VkPhysicalDeviceVideoEncodeRgbConversionFeaturesVALVE {
pub mut:
	sType                    StructureType = StructureType.physical_device_video_encode_rgb_conversion_features_valve
	pNext                    voidptr       = unsafe { nil }
	videoEncodeRgbConversion Bool32
}

// VideoEncodeRgbConversionCapabilitiesVALVE extends VkVideoCapabilitiesKHR
pub type VideoEncodeRgbConversionCapabilitiesVALVE = C.VkVideoEncodeRgbConversionCapabilitiesVALVE

@[typedef]
pub struct C.VkVideoEncodeRgbConversionCapabilitiesVALVE {
pub mut:
	sType          StructureType = StructureType.video_encode_rgb_conversion_capabilities_valve
	pNext          voidptr       = unsafe { nil }
	rgbModels      VideoEncodeRgbModelConversionFlagsVALVE
	rgbRanges      VideoEncodeRgbRangeCompressionFlagsVALVE
	xChromaOffsets VideoEncodeRgbChromaOffsetFlagsVALVE
	yChromaOffsets VideoEncodeRgbChromaOffsetFlagsVALVE
}

// VideoEncodeProfileRgbConversionInfoVALVE extends VkVideoProfileInfoKHR
pub type VideoEncodeProfileRgbConversionInfoVALVE = C.VkVideoEncodeProfileRgbConversionInfoVALVE

@[typedef]
pub struct C.VkVideoEncodeProfileRgbConversionInfoVALVE {
pub mut:
	sType                      StructureType = StructureType.video_encode_profile_rgb_conversion_info_valve
	pNext                      voidptr       = unsafe { nil }
	performEncodeRgbConversion Bool32
}

// VideoEncodeSessionRgbConversionCreateInfoVALVE extends VkVideoSessionCreateInfoKHR
pub type VideoEncodeSessionRgbConversionCreateInfoVALVE = C.VkVideoEncodeSessionRgbConversionCreateInfoVALVE

@[typedef]
pub struct C.VkVideoEncodeSessionRgbConversionCreateInfoVALVE {
pub mut:
	sType         StructureType = StructureType.video_encode_session_rgb_conversion_create_info_valve
	pNext         voidptr       = unsafe { nil }
	rgbModel      VideoEncodeRgbModelConversionFlagBitsVALVE
	rgbRange      VideoEncodeRgbRangeCompressionFlagBitsVALVE
	xChromaOffset VideoEncodeRgbChromaOffsetFlagBitsVALVE
	yChromaOffset VideoEncodeRgbChromaOffsetFlagBitsVALVE
}

pub const ext_image_view_min_lod_spec_version = 1
pub const ext_image_view_min_lod_extension_name = c'VK_EXT_image_view_min_lod'
// PhysicalDeviceImageViewMinLodFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceImageViewMinLodFeaturesEXT = C.VkPhysicalDeviceImageViewMinLodFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceImageViewMinLodFeaturesEXT {
pub mut:
	sType  StructureType = StructureType.physical_device_image_view_min_lod_features_ext
	pNext  voidptr       = unsafe { nil }
	minLod Bool32
}

// ImageViewMinLodCreateInfoEXT extends VkImageViewCreateInfo
pub type ImageViewMinLodCreateInfoEXT = C.VkImageViewMinLodCreateInfoEXT

@[typedef]
pub struct C.VkImageViewMinLodCreateInfoEXT {
pub mut:
	sType  StructureType = StructureType.image_view_min_lod_create_info_ext
	pNext  voidptr       = unsafe { nil }
	minLod f32
}

pub const ext_multi_draw_spec_version = 1
pub const ext_multi_draw_extension_name = c'VK_EXT_multi_draw'
// PhysicalDeviceMultiDrawFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMultiDrawFeaturesEXT = C.VkPhysicalDeviceMultiDrawFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMultiDrawFeaturesEXT {
pub mut:
	sType     StructureType = StructureType.physical_device_multi_draw_features_ext
	pNext     voidptr       = unsafe { nil }
	multiDraw Bool32
}

// PhysicalDeviceMultiDrawPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMultiDrawPropertiesEXT = C.VkPhysicalDeviceMultiDrawPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMultiDrawPropertiesEXT {
pub mut:
	sType             StructureType = StructureType.physical_device_multi_draw_properties_ext
	pNext             voidptr       = unsafe { nil }
	maxMultiDrawCount u32
}

pub type MultiDrawInfoEXT = C.VkMultiDrawInfoEXT

@[typedef]
pub struct C.VkMultiDrawInfoEXT {
pub mut:
	firstVertex u32
	vertexCount u32
}

pub type MultiDrawIndexedInfoEXT = C.VkMultiDrawIndexedInfoEXT

@[typedef]
pub struct C.VkMultiDrawIndexedInfoEXT {
pub mut:
	firstIndex   u32
	indexCount   u32
	vertexOffset i32
}

@[keep_args_alive]
fn C.vkCmdDrawMultiEXT(command_buffer CommandBuffer, draw_count u32, p_vertex_info &MultiDrawInfoEXT, instance_count u32, first_instance u32, stride u32)

pub type PFN_vkCmdDrawMultiEXT = fn (command_buffer CommandBuffer, draw_count u32, p_vertex_info &MultiDrawInfoEXT, instance_count u32, first_instance u32, stride u32)

@[inline]
pub fn cmd_draw_multi_ext(command_buffer CommandBuffer,
	draw_count u32,
	p_vertex_info &MultiDrawInfoEXT,
	instance_count u32,
	first_instance u32,
	stride u32) {
	C.vkCmdDrawMultiEXT(command_buffer, draw_count, p_vertex_info, instance_count, first_instance,
		stride)
}

@[keep_args_alive]
fn C.vkCmdDrawMultiIndexedEXT(command_buffer CommandBuffer, draw_count u32, p_index_info &MultiDrawIndexedInfoEXT, instance_count u32, first_instance u32, stride u32, p_vertex_offset &i32)

pub type PFN_vkCmdDrawMultiIndexedEXT = fn (command_buffer CommandBuffer, draw_count u32, p_index_info &MultiDrawIndexedInfoEXT, instance_count u32, first_instance u32, stride u32, p_vertex_offset &i32)

@[inline]
pub fn cmd_draw_multi_indexed_ext(command_buffer CommandBuffer,
	draw_count u32,
	p_index_info &MultiDrawIndexedInfoEXT,
	instance_count u32,
	first_instance u32,
	stride u32,
	p_vertex_offset &i32) {
	C.vkCmdDrawMultiIndexedEXT(command_buffer, draw_count, p_index_info, instance_count,
		first_instance, stride, p_vertex_offset)
}

pub const ext_image_2d_view_of_3d_spec_version = 1
pub const ext_image_2d_view_of_3d_extension_name = c'VK_EXT_image_2d_view_of_3d'
// PhysicalDeviceImage2DViewOf3DFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceImage2DViewOf3DFeaturesEXT = C.VkPhysicalDeviceImage2DViewOf3DFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceImage2DViewOf3DFeaturesEXT {
pub mut:
	sType             StructureType = StructureType.physical_device_image2d_view_of3d_features_ext
	pNext             voidptr       = unsafe { nil }
	image2DViewOf3D   Bool32
	sampler2DViewOf3D Bool32
}

pub const ext_shader_tile_image_spec_version = 1
pub const ext_shader_tile_image_extension_name = c'VK_EXT_shader_tile_image'
// PhysicalDeviceShaderTileImageFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderTileImageFeaturesEXT = C.VkPhysicalDeviceShaderTileImageFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderTileImageFeaturesEXT {
pub mut:
	sType                            StructureType = StructureType.physical_device_shader_tile_image_features_ext
	pNext                            voidptr       = unsafe { nil }
	shaderTileImageColorReadAccess   Bool32
	shaderTileImageDepthReadAccess   Bool32
	shaderTileImageStencilReadAccess Bool32
}

// PhysicalDeviceShaderTileImagePropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceShaderTileImagePropertiesEXT = C.VkPhysicalDeviceShaderTileImagePropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderTileImagePropertiesEXT {
pub mut:
	sType                                            StructureType = StructureType.physical_device_shader_tile_image_properties_ext
	pNext                                            voidptr       = unsafe { nil }
	shaderTileImageCoherentReadAccelerated           Bool32
	shaderTileImageReadSampleFromPixelRateInvocation Bool32
	shaderTileImageReadFromHelperInvocation          Bool32
}

// Pointer to VkMicromapEXT_T
pub type MicromapEXT = voidptr

pub const ext_opacity_micromap_spec_version = 2
pub const ext_opacity_micromap_extension_name = c'VK_EXT_opacity_micromap'

pub enum MicromapTypeEXT as u32 {
	opacity_micromap = 0
	max_enum_ext     = max_int
}

pub enum BuildMicromapModeEXT as u32 {
	build        = 0
	max_enum_ext = max_int
}

pub enum CopyMicromapModeEXT as u32 {
	clone        = 0
	serialize    = 1
	deserialize  = 2
	compact      = 3
	max_enum_ext = max_int
}

pub enum OpacityMicromapFormatEXT as u32 {
	_2_state     = 1
	_4_state     = 2
	max_enum_ext = max_int
}

pub enum OpacityMicromapSpecialIndexEXT {
	fully_transparent                            = -1
	fully_opaque                                 = -2
	fully_unknown_transparent                    = -3
	fully_unknown_opaque                         = -4
	cluster_geometry_disable_opacity_micromap_nv = -5
	max_enum_ext                                 = max_int
}

pub enum AccelerationStructureCompatibilityKHR as u32 {
	compatible   = 0
	incompatible = 1
	max_enum_khr = max_int
}

pub enum AccelerationStructureBuildTypeKHR as u32 {
	host           = 0
	device         = 1
	host_or_device = 2
	max_enum_khr   = max_int
}

pub enum BuildMicromapFlagBitsEXT as u32 {
	prefer_fast_trace = u32(0x00000001)
	prefer_fast_build = u32(0x00000002)
	allow_compaction  = u32(0x00000004)
	max_enum_ext      = max_int
}
pub type BuildMicromapFlagsEXT = u32

pub enum MicromapCreateFlagBitsEXT as u32 {
	device_address_capture_replay = u32(0x00000001)
	max_enum_ext                  = max_int
}
pub type MicromapCreateFlagsEXT = u32
pub type MicromapUsageEXT = C.VkMicromapUsageEXT

@[typedef]
pub struct C.VkMicromapUsageEXT {
pub mut:
	count            u32
	subdivisionLevel u32
	format           u32
}

pub type DeviceOrHostAddressKHR = C.VkDeviceOrHostAddressKHR

@[typedef]
pub union C.VkDeviceOrHostAddressKHR {
pub mut:
	deviceAddress DeviceAddress
	hostAddress   voidptr
}

pub type MicromapBuildInfoEXT = C.VkMicromapBuildInfoEXT

@[typedef]
pub struct C.VkMicromapBuildInfoEXT {
pub mut:
	sType               StructureType = StructureType.micromap_build_info_ext
	pNext               voidptr       = unsafe { nil }
	type                MicromapTypeEXT
	flags               BuildMicromapFlagsEXT
	mode                BuildMicromapModeEXT
	dstMicromap         MicromapEXT
	usageCountsCount    u32
	pUsageCounts        &MicromapUsageEXT
	ppUsageCounts       &&MicromapUsageEXT
	data                DeviceOrHostAddressConstKHR
	scratchData         DeviceOrHostAddressKHR
	triangleArray       DeviceOrHostAddressConstKHR
	triangleArrayStride DeviceSize
}

pub type MicromapCreateInfoEXT = C.VkMicromapCreateInfoEXT

@[typedef]
pub struct C.VkMicromapCreateInfoEXT {
pub mut:
	sType         StructureType = StructureType.micromap_create_info_ext
	pNext         voidptr       = unsafe { nil }
	createFlags   MicromapCreateFlagsEXT
	buffer        Buffer
	offset        DeviceSize
	size          DeviceSize
	type          MicromapTypeEXT
	deviceAddress DeviceAddress
}

// PhysicalDeviceOpacityMicromapFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceOpacityMicromapFeaturesEXT = C.VkPhysicalDeviceOpacityMicromapFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceOpacityMicromapFeaturesEXT {
pub mut:
	sType                 StructureType = StructureType.physical_device_opacity_micromap_features_ext
	pNext                 voidptr       = unsafe { nil }
	micromap              Bool32
	micromapCaptureReplay Bool32
	micromapHostCommands  Bool32
}

// PhysicalDeviceOpacityMicromapPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceOpacityMicromapPropertiesEXT = C.VkPhysicalDeviceOpacityMicromapPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceOpacityMicromapPropertiesEXT {
pub mut:
	sType                            StructureType = StructureType.physical_device_opacity_micromap_properties_ext
	pNext                            voidptr       = unsafe { nil }
	maxOpacity2StateSubdivisionLevel u32
	maxOpacity4StateSubdivisionLevel u32
}

pub type MicromapVersionInfoEXT = C.VkMicromapVersionInfoEXT

@[typedef]
pub struct C.VkMicromapVersionInfoEXT {
pub mut:
	sType        StructureType = StructureType.micromap_version_info_ext
	pNext        voidptr       = unsafe { nil }
	pVersionData &u8
}

pub type CopyMicromapToMemoryInfoEXT = C.VkCopyMicromapToMemoryInfoEXT

@[typedef]
pub struct C.VkCopyMicromapToMemoryInfoEXT {
pub mut:
	sType StructureType = StructureType.copy_micromap_to_memory_info_ext
	pNext voidptr       = unsafe { nil }
	src   MicromapEXT
	dst   DeviceOrHostAddressKHR
	mode  CopyMicromapModeEXT
}

pub type CopyMemoryToMicromapInfoEXT = C.VkCopyMemoryToMicromapInfoEXT

@[typedef]
pub struct C.VkCopyMemoryToMicromapInfoEXT {
pub mut:
	sType StructureType = StructureType.copy_memory_to_micromap_info_ext
	pNext voidptr       = unsafe { nil }
	src   DeviceOrHostAddressConstKHR
	dst   MicromapEXT
	mode  CopyMicromapModeEXT
}

pub type CopyMicromapInfoEXT = C.VkCopyMicromapInfoEXT

@[typedef]
pub struct C.VkCopyMicromapInfoEXT {
pub mut:
	sType StructureType = StructureType.copy_micromap_info_ext
	pNext voidptr       = unsafe { nil }
	src   MicromapEXT
	dst   MicromapEXT
	mode  CopyMicromapModeEXT
}

pub type MicromapBuildSizesInfoEXT = C.VkMicromapBuildSizesInfoEXT

@[typedef]
pub struct C.VkMicromapBuildSizesInfoEXT {
pub mut:
	sType            StructureType = StructureType.micromap_build_sizes_info_ext
	pNext            voidptr       = unsafe { nil }
	micromapSize     DeviceSize
	buildScratchSize DeviceSize
	discardable      Bool32
}

// AccelerationStructureTrianglesOpacityMicromapEXT extends VkAccelerationStructureGeometryTrianglesDataKHR,VkAccelerationStructureDenseGeometryFormatTrianglesDataAMDX
pub type AccelerationStructureTrianglesOpacityMicromapEXT = C.VkAccelerationStructureTrianglesOpacityMicromapEXT

@[typedef]
pub struct C.VkAccelerationStructureTrianglesOpacityMicromapEXT {
pub mut:
	sType            StructureType = StructureType.acceleration_structure_triangles_opacity_micromap_ext
	pNext            voidptr       = unsafe { nil }
	indexType        IndexType
	indexBuffer      DeviceOrHostAddressConstKHR
	indexStride      DeviceSize
	baseTriangle     u32
	usageCountsCount u32
	pUsageCounts     &MicromapUsageEXT
	ppUsageCounts    &&MicromapUsageEXT
	micromap         MicromapEXT
}

pub type MicromapTriangleEXT = C.VkMicromapTriangleEXT

@[typedef]
pub struct C.VkMicromapTriangleEXT {
pub mut:
	dataOffset       u32
	subdivisionLevel u16
	format           u16
}

@[keep_args_alive]
fn C.vkCreateMicromapEXT(device Device, p_create_info &MicromapCreateInfoEXT, p_allocator &AllocationCallbacks, p_micromap &MicromapEXT) Result

pub type PFN_vkCreateMicromapEXT = fn (device Device, p_create_info &MicromapCreateInfoEXT, p_allocator &AllocationCallbacks, p_micromap &MicromapEXT) Result

@[inline]
pub fn create_micromap_ext(device Device,
	p_create_info &MicromapCreateInfoEXT,
	p_allocator &AllocationCallbacks,
	p_micromap &MicromapEXT) Result {
	return C.vkCreateMicromapEXT(device, p_create_info, p_allocator, p_micromap)
}

@[keep_args_alive]
fn C.vkDestroyMicromapEXT(device Device, micromap MicromapEXT, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyMicromapEXT = fn (device Device, micromap MicromapEXT, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_micromap_ext(device Device,
	micromap MicromapEXT,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyMicromapEXT(device, micromap, p_allocator)
}

@[keep_args_alive]
fn C.vkCmdBuildMicromapsEXT(command_buffer CommandBuffer, info_count u32, p_infos &MicromapBuildInfoEXT)

pub type PFN_vkCmdBuildMicromapsEXT = fn (command_buffer CommandBuffer, info_count u32, p_infos &MicromapBuildInfoEXT)

@[inline]
pub fn cmd_build_micromaps_ext(command_buffer CommandBuffer,
	info_count u32,
	p_infos &MicromapBuildInfoEXT) {
	C.vkCmdBuildMicromapsEXT(command_buffer, info_count, p_infos)
}

@[keep_args_alive]
fn C.vkBuildMicromapsEXT(device Device, deferred_operation DeferredOperationKHR, info_count u32, p_infos &MicromapBuildInfoEXT) Result

pub type PFN_vkBuildMicromapsEXT = fn (device Device, deferred_operation DeferredOperationKHR, info_count u32, p_infos &MicromapBuildInfoEXT) Result

@[inline]
pub fn build_micromaps_ext(device Device,
	deferred_operation DeferredOperationKHR,
	info_count u32,
	p_infos &MicromapBuildInfoEXT) Result {
	return C.vkBuildMicromapsEXT(device, deferred_operation, info_count, p_infos)
}

@[keep_args_alive]
fn C.vkCopyMicromapEXT(device Device, deferred_operation DeferredOperationKHR, p_info &CopyMicromapInfoEXT) Result

pub type PFN_vkCopyMicromapEXT = fn (device Device, deferred_operation DeferredOperationKHR, p_info &CopyMicromapInfoEXT) Result

@[inline]
pub fn copy_micromap_ext(device Device,
	deferred_operation DeferredOperationKHR,
	p_info &CopyMicromapInfoEXT) Result {
	return C.vkCopyMicromapEXT(device, deferred_operation, p_info)
}

@[keep_args_alive]
fn C.vkCopyMicromapToMemoryEXT(device Device, deferred_operation DeferredOperationKHR, p_info &CopyMicromapToMemoryInfoEXT) Result

pub type PFN_vkCopyMicromapToMemoryEXT = fn (device Device, deferred_operation DeferredOperationKHR, p_info &CopyMicromapToMemoryInfoEXT) Result

@[inline]
pub fn copy_micromap_to_memory_ext(device Device,
	deferred_operation DeferredOperationKHR,
	p_info &CopyMicromapToMemoryInfoEXT) Result {
	return C.vkCopyMicromapToMemoryEXT(device, deferred_operation, p_info)
}

@[keep_args_alive]
fn C.vkCopyMemoryToMicromapEXT(device Device, deferred_operation DeferredOperationKHR, p_info &CopyMemoryToMicromapInfoEXT) Result

pub type PFN_vkCopyMemoryToMicromapEXT = fn (device Device, deferred_operation DeferredOperationKHR, p_info &CopyMemoryToMicromapInfoEXT) Result

@[inline]
pub fn copy_memory_to_micromap_ext(device Device,
	deferred_operation DeferredOperationKHR,
	p_info &CopyMemoryToMicromapInfoEXT) Result {
	return C.vkCopyMemoryToMicromapEXT(device, deferred_operation, p_info)
}

@[keep_args_alive]
fn C.vkWriteMicromapsPropertiesEXT(device Device, micromap_count u32, p_micromaps &MicromapEXT, query_type QueryType, data_size usize, p_data voidptr, stride usize) Result

pub type PFN_vkWriteMicromapsPropertiesEXT = fn (device Device, micromap_count u32, p_micromaps &MicromapEXT, query_type QueryType, data_size usize, p_data voidptr, stride usize) Result

@[inline]
pub fn write_micromaps_properties_ext(device Device,
	micromap_count u32,
	p_micromaps &MicromapEXT,
	query_type QueryType,
	data_size usize,
	p_data voidptr,
	stride usize) Result {
	return C.vkWriteMicromapsPropertiesEXT(device, micromap_count, p_micromaps, query_type,
		data_size, p_data, stride)
}

@[keep_args_alive]
fn C.vkCmdCopyMicromapEXT(command_buffer CommandBuffer, p_info &CopyMicromapInfoEXT)

pub type PFN_vkCmdCopyMicromapEXT = fn (command_buffer CommandBuffer, p_info &CopyMicromapInfoEXT)

@[inline]
pub fn cmd_copy_micromap_ext(command_buffer CommandBuffer,
	p_info &CopyMicromapInfoEXT) {
	C.vkCmdCopyMicromapEXT(command_buffer, p_info)
}

@[keep_args_alive]
fn C.vkCmdCopyMicromapToMemoryEXT(command_buffer CommandBuffer, p_info &CopyMicromapToMemoryInfoEXT)

pub type PFN_vkCmdCopyMicromapToMemoryEXT = fn (command_buffer CommandBuffer, p_info &CopyMicromapToMemoryInfoEXT)

@[inline]
pub fn cmd_copy_micromap_to_memory_ext(command_buffer CommandBuffer,
	p_info &CopyMicromapToMemoryInfoEXT) {
	C.vkCmdCopyMicromapToMemoryEXT(command_buffer, p_info)
}

@[keep_args_alive]
fn C.vkCmdCopyMemoryToMicromapEXT(command_buffer CommandBuffer, p_info &CopyMemoryToMicromapInfoEXT)

pub type PFN_vkCmdCopyMemoryToMicromapEXT = fn (command_buffer CommandBuffer, p_info &CopyMemoryToMicromapInfoEXT)

@[inline]
pub fn cmd_copy_memory_to_micromap_ext(command_buffer CommandBuffer,
	p_info &CopyMemoryToMicromapInfoEXT) {
	C.vkCmdCopyMemoryToMicromapEXT(command_buffer, p_info)
}

@[keep_args_alive]
fn C.vkCmdWriteMicromapsPropertiesEXT(command_buffer CommandBuffer, micromap_count u32, p_micromaps &MicromapEXT, query_type QueryType, query_pool QueryPool, first_query u32)

pub type PFN_vkCmdWriteMicromapsPropertiesEXT = fn (command_buffer CommandBuffer, micromap_count u32, p_micromaps &MicromapEXT, query_type QueryType, query_pool QueryPool, first_query u32)

@[inline]
pub fn cmd_write_micromaps_properties_ext(command_buffer CommandBuffer,
	micromap_count u32,
	p_micromaps &MicromapEXT,
	query_type QueryType,
	query_pool QueryPool,
	first_query u32) {
	C.vkCmdWriteMicromapsPropertiesEXT(command_buffer, micromap_count, p_micromaps, query_type,
		query_pool, first_query)
}

@[keep_args_alive]
fn C.vkGetDeviceMicromapCompatibilityEXT(device Device, p_version_info &MicromapVersionInfoEXT, p_compatibility &AccelerationStructureCompatibilityKHR)

pub type PFN_vkGetDeviceMicromapCompatibilityEXT = fn (device Device, p_version_info &MicromapVersionInfoEXT, p_compatibility &AccelerationStructureCompatibilityKHR)

@[inline]
pub fn get_device_micromap_compatibility_ext(device Device,
	p_version_info &MicromapVersionInfoEXT,
	p_compatibility &AccelerationStructureCompatibilityKHR) {
	C.vkGetDeviceMicromapCompatibilityEXT(device, p_version_info, p_compatibility)
}

@[keep_args_alive]
fn C.vkGetMicromapBuildSizesEXT(device Device, build_type AccelerationStructureBuildTypeKHR, p_build_info &MicromapBuildInfoEXT, mut p_size_info MicromapBuildSizesInfoEXT)

pub type PFN_vkGetMicromapBuildSizesEXT = fn (device Device, build_type AccelerationStructureBuildTypeKHR, p_build_info &MicromapBuildInfoEXT, mut p_size_info MicromapBuildSizesInfoEXT)

@[inline]
pub fn get_micromap_build_sizes_ext(device Device,
	build_type AccelerationStructureBuildTypeKHR,
	p_build_info &MicromapBuildInfoEXT,
	mut p_size_info MicromapBuildSizesInfoEXT) {
	C.vkGetMicromapBuildSizesEXT(device, build_type, p_build_info, mut p_size_info)
}

pub const ext_load_store_op_none_spec_version = 1
pub const ext_load_store_op_none_extension_name = c'VK_EXT_load_store_op_none'

pub const huawei_cluster_culling_shader_spec_version = 3
pub const huawei_cluster_culling_shader_extension_name = c'VK_HAWEI_cluster_culling_shader'
// PhysicalDeviceClusterCullingShaderFeaturesHUAWEI extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceClusterCullingShaderFeaturesHUAWEI = C.VkPhysicalDeviceClusterCullingShaderFeaturesHUAWEI

@[typedef]
pub struct C.VkPhysicalDeviceClusterCullingShaderFeaturesHUAWEI {
pub mut:
	sType                         StructureType = StructureType.physical_device_cluster_culling_shader_features_huawei
	pNext                         voidptr       = unsafe { nil }
	clustercullingShader          Bool32
	multiviewClusterCullingShader Bool32
}

// PhysicalDeviceClusterCullingShaderPropertiesHUAWEI extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceClusterCullingShaderPropertiesHUAWEI = C.VkPhysicalDeviceClusterCullingShaderPropertiesHUAWEI

@[typedef]
pub struct C.VkPhysicalDeviceClusterCullingShaderPropertiesHUAWEI {
pub mut:
	sType                         StructureType = StructureType.physical_device_cluster_culling_shader_properties_huawei
	pNext                         voidptr       = unsafe { nil }
	maxWorkGroupCount             [3]u32
	maxWorkGroupSize              [3]u32
	maxOutputClusterCount         u32
	indirectBufferOffsetAlignment DeviceSize
}

// PhysicalDeviceClusterCullingShaderVrsFeaturesHUAWEI extends VkPhysicalDeviceClusterCullingShaderFeaturesHUAWEI
pub type PhysicalDeviceClusterCullingShaderVrsFeaturesHUAWEI = C.VkPhysicalDeviceClusterCullingShaderVrsFeaturesHUAWEI

@[typedef]
pub struct C.VkPhysicalDeviceClusterCullingShaderVrsFeaturesHUAWEI {
pub mut:
	sType              StructureType = StructureType.physical_device_cluster_culling_shader_vrs_features_huawei
	pNext              voidptr       = unsafe { nil }
	clusterShadingRate Bool32
}

@[keep_args_alive]
fn C.vkCmdDrawClusterHUAWEI(command_buffer CommandBuffer, group_count_x u32, group_count_y u32, group_count_z u32)

pub type PFN_vkCmdDrawClusterHUAWEI = fn (command_buffer CommandBuffer, group_count_x u32, group_count_y u32, group_count_z u32)

@[inline]
pub fn cmd_draw_cluster_huawei(command_buffer CommandBuffer,
	group_count_x u32,
	group_count_y u32,
	group_count_z u32) {
	C.vkCmdDrawClusterHUAWEI(command_buffer, group_count_x, group_count_y, group_count_z)
}

@[keep_args_alive]
fn C.vkCmdDrawClusterIndirectHUAWEI(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize)

pub type PFN_vkCmdDrawClusterIndirectHUAWEI = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize)

@[inline]
pub fn cmd_draw_cluster_indirect_huawei(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize) {
	C.vkCmdDrawClusterIndirectHUAWEI(command_buffer, buffer, offset)
}

pub const ext_border_color_swizzle_spec_version = 1
pub const ext_border_color_swizzle_extension_name = c'VK_EXT_border_color_swizzle'
// PhysicalDeviceBorderColorSwizzleFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceBorderColorSwizzleFeaturesEXT = C.VkPhysicalDeviceBorderColorSwizzleFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceBorderColorSwizzleFeaturesEXT {
pub mut:
	sType                       StructureType = StructureType.physical_device_border_color_swizzle_features_ext
	pNext                       voidptr       = unsafe { nil }
	borderColorSwizzle          Bool32
	borderColorSwizzleFromImage Bool32
}

// SamplerBorderColorComponentMappingCreateInfoEXT extends VkSamplerCreateInfo
pub type SamplerBorderColorComponentMappingCreateInfoEXT = C.VkSamplerBorderColorComponentMappingCreateInfoEXT

@[typedef]
pub struct C.VkSamplerBorderColorComponentMappingCreateInfoEXT {
pub mut:
	sType      StructureType = StructureType.sampler_border_color_component_mapping_create_info_ext
	pNext      voidptr       = unsafe { nil }
	components ComponentMapping
	srgb       Bool32
}

pub const ext_pageable_device_local_memory_spec_version = 1
pub const ext_pageable_device_local_memory_extension_name = c'VK_EXT_pageable_device_local_memory'
// PhysicalDevicePageableDeviceLocalMemoryFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePageableDeviceLocalMemoryFeaturesEXT = C.VkPhysicalDevicePageableDeviceLocalMemoryFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDevicePageableDeviceLocalMemoryFeaturesEXT {
pub mut:
	sType                     StructureType = StructureType.physical_device_pageable_device_local_memory_features_ext
	pNext                     voidptr       = unsafe { nil }
	pageableDeviceLocalMemory Bool32
}

@[keep_args_alive]
fn C.vkSetDeviceMemoryPriorityEXT(device Device, memory DeviceMemory, priority f32)

pub type PFN_vkSetDeviceMemoryPriorityEXT = fn (device Device, memory DeviceMemory, priority f32)

@[inline]
pub fn set_device_memory_priority_ext(device Device,
	memory DeviceMemory,
	priority f32) {
	C.vkSetDeviceMemoryPriorityEXT(device, memory, priority)
}

pub const arm_shader_core_properties_spec_version = 1
pub const arm_shader_core_properties_extension_name = c'VK_ARM_shader_core_properties'
// PhysicalDeviceShaderCorePropertiesARM extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceShaderCorePropertiesARM = C.VkPhysicalDeviceShaderCorePropertiesARM

@[typedef]
pub struct C.VkPhysicalDeviceShaderCorePropertiesARM {
pub mut:
	sType     StructureType = StructureType.physical_device_shader_core_properties_arm
	pNext     voidptr       = unsafe { nil }
	pixelRate u32
	texelRate u32
	fmaRate   u32
}

pub const arm_scheduling_controls_spec_version = 1
pub const arm_scheduling_controls_extension_name = c'VK_ARM_scheduling_controls'

pub type PhysicalDeviceSchedulingControlsFlagsARM = u64

// Flag bits for PhysicalDeviceSchedulingControlsFlagBitsARM
pub type PhysicalDeviceSchedulingControlsFlagBitsARM = u64

pub const physical_device_scheduling_controls_shader_core_count_arm = u64(0x00000001)

// DeviceQueueShaderCoreControlCreateInfoARM extends VkDeviceQueueCreateInfo,VkDeviceCreateInfo
pub type DeviceQueueShaderCoreControlCreateInfoARM = C.VkDeviceQueueShaderCoreControlCreateInfoARM

@[typedef]
pub struct C.VkDeviceQueueShaderCoreControlCreateInfoARM {
pub mut:
	sType           StructureType = StructureType.device_queue_shader_core_control_create_info_arm
	pNext           voidptr       = unsafe { nil }
	shaderCoreCount u32
}

// PhysicalDeviceSchedulingControlsFeaturesARM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceSchedulingControlsFeaturesARM = C.VkPhysicalDeviceSchedulingControlsFeaturesARM

@[typedef]
pub struct C.VkPhysicalDeviceSchedulingControlsFeaturesARM {
pub mut:
	sType              StructureType = StructureType.physical_device_scheduling_controls_features_arm
	pNext              voidptr       = unsafe { nil }
	schedulingControls Bool32
}

// PhysicalDeviceSchedulingControlsPropertiesARM extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceSchedulingControlsPropertiesARM = C.VkPhysicalDeviceSchedulingControlsPropertiesARM

@[typedef]
pub struct C.VkPhysicalDeviceSchedulingControlsPropertiesARM {
pub mut:
	sType                   StructureType = StructureType.physical_device_scheduling_controls_properties_arm
	pNext                   voidptr       = unsafe { nil }
	schedulingControlsFlags PhysicalDeviceSchedulingControlsFlagsARM
}

pub const ext_image_sliced_view_of_3d_spec_version = 1
pub const ext_image_sliced_view_of_3d_extension_name = c'VK_EXT_image_sliced_view_of_3d'
pub const remaining_3d_slices_ext = ~u32(0)
// PhysicalDeviceImageSlicedViewOf3DFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceImageSlicedViewOf3DFeaturesEXT = C.VkPhysicalDeviceImageSlicedViewOf3DFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceImageSlicedViewOf3DFeaturesEXT {
pub mut:
	sType               StructureType = StructureType.physical_device_image_sliced_view_of3d_features_ext
	pNext               voidptr       = unsafe { nil }
	imageSlicedViewOf3D Bool32
}

// ImageViewSlicedCreateInfoEXT extends VkImageViewCreateInfo
pub type ImageViewSlicedCreateInfoEXT = C.VkImageViewSlicedCreateInfoEXT

@[typedef]
pub struct C.VkImageViewSlicedCreateInfoEXT {
pub mut:
	sType       StructureType = StructureType.image_view_sliced_create_info_ext
	pNext       voidptr       = unsafe { nil }
	sliceOffset u32
	sliceCount  u32
}

pub const valve_descriptor_set_host_mapping_spec_version = 1
pub const valve_descriptor_set_host_mapping_extension_name = c'VK_VAVE_descriptor_set_host_mapping'
// PhysicalDeviceDescriptorSetHostMappingFeaturesVALVE extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDescriptorSetHostMappingFeaturesVALVE = C.VkPhysicalDeviceDescriptorSetHostMappingFeaturesVALVE

@[typedef]
pub struct C.VkPhysicalDeviceDescriptorSetHostMappingFeaturesVALVE {
pub mut:
	sType                    StructureType = StructureType.physical_device_descriptor_set_host_mapping_features_valve
	pNext                    voidptr       = unsafe { nil }
	descriptorSetHostMapping Bool32
}

pub type DescriptorSetBindingReferenceVALVE = C.VkDescriptorSetBindingReferenceVALVE

@[typedef]
pub struct C.VkDescriptorSetBindingReferenceVALVE {
pub mut:
	sType               StructureType = StructureType.descriptor_set_binding_reference_valve
	pNext               voidptr       = unsafe { nil }
	descriptorSetLayout DescriptorSetLayout
	binding             u32
}

pub type DescriptorSetLayoutHostMappingInfoVALVE = C.VkDescriptorSetLayoutHostMappingInfoVALVE

@[typedef]
pub struct C.VkDescriptorSetLayoutHostMappingInfoVALVE {
pub mut:
	sType            StructureType = StructureType.descriptor_set_layout_host_mapping_info_valve
	pNext            voidptr       = unsafe { nil }
	descriptorOffset usize
	descriptorSize   u32
}

@[keep_args_alive]
fn C.vkGetDescriptorSetLayoutHostMappingInfoVALVE(device Device, p_binding_reference &DescriptorSetBindingReferenceVALVE, mut p_host_mapping DescriptorSetLayoutHostMappingInfoVALVE)

pub type PFN_vkGetDescriptorSetLayoutHostMappingInfoVALVE = fn (device Device, p_binding_reference &DescriptorSetBindingReferenceVALVE, mut p_host_mapping DescriptorSetLayoutHostMappingInfoVALVE)

@[inline]
pub fn get_descriptor_set_layout_host_mapping_info_valve(device Device,
	p_binding_reference &DescriptorSetBindingReferenceVALVE,
	mut p_host_mapping DescriptorSetLayoutHostMappingInfoVALVE) {
	C.vkGetDescriptorSetLayoutHostMappingInfoVALVE(device, p_binding_reference, mut p_host_mapping)
}

@[keep_args_alive]
fn C.vkGetDescriptorSetHostMappingVALVE(device Device, descriptor_set DescriptorSet, pp_data &voidptr)

pub type PFN_vkGetDescriptorSetHostMappingVALVE = fn (device Device, descriptor_set DescriptorSet, pp_data &voidptr)

@[inline]
pub fn get_descriptor_set_host_mapping_valve(device Device,
	descriptor_set DescriptorSet,
	pp_data &voidptr) {
	C.vkGetDescriptorSetHostMappingVALVE(device, descriptor_set, pp_data)
}

pub const ext_depth_clamp_zero_one_spec_version = 1
pub const ext_depth_clamp_zero_one_extension_name = c'VK_EXT_depth_clamp_zero_one'

pub type PhysicalDeviceDepthClampZeroOneFeaturesEXT = C.VkPhysicalDeviceDepthClampZeroOneFeaturesKHR

pub const ext_non_seamless_cube_map_spec_version = 1
pub const ext_non_seamless_cube_map_extension_name = c'VK_EXT_non_seamless_cube_map'
// PhysicalDeviceNonSeamlessCubeMapFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceNonSeamlessCubeMapFeaturesEXT = C.VkPhysicalDeviceNonSeamlessCubeMapFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceNonSeamlessCubeMapFeaturesEXT {
pub mut:
	sType              StructureType = StructureType.physical_device_non_seamless_cube_map_features_ext
	pNext              voidptr       = unsafe { nil }
	nonSeamlessCubeMap Bool32
}

pub const arm_render_pass_striped_spec_version = 1
pub const arm_render_pass_striped_extension_name = c'VK_ARM_render_pass_striped'
// PhysicalDeviceRenderPassStripedFeaturesARM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRenderPassStripedFeaturesARM = C.VkPhysicalDeviceRenderPassStripedFeaturesARM

@[typedef]
pub struct C.VkPhysicalDeviceRenderPassStripedFeaturesARM {
pub mut:
	sType             StructureType = StructureType.physical_device_render_pass_striped_features_arm
	pNext             voidptr       = unsafe { nil }
	renderPassStriped Bool32
}

// PhysicalDeviceRenderPassStripedPropertiesARM extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceRenderPassStripedPropertiesARM = C.VkPhysicalDeviceRenderPassStripedPropertiesARM

@[typedef]
pub struct C.VkPhysicalDeviceRenderPassStripedPropertiesARM {
pub mut:
	sType                       StructureType = StructureType.physical_device_render_pass_striped_properties_arm
	pNext                       voidptr       = unsafe { nil }
	renderPassStripeGranularity Extent2D
	maxRenderPassStripes        u32
}

pub type RenderPassStripeInfoARM = C.VkRenderPassStripeInfoARM

@[typedef]
pub struct C.VkRenderPassStripeInfoARM {
pub mut:
	sType      StructureType = StructureType.render_pass_stripe_info_arm
	pNext      voidptr       = unsafe { nil }
	stripeArea Rect2D
}

// RenderPassStripeBeginInfoARM extends VkRenderingInfo,VkRenderPassBeginInfo
pub type RenderPassStripeBeginInfoARM = C.VkRenderPassStripeBeginInfoARM

@[typedef]
pub struct C.VkRenderPassStripeBeginInfoARM {
pub mut:
	sType           StructureType = StructureType.render_pass_stripe_begin_info_arm
	pNext           voidptr       = unsafe { nil }
	stripeInfoCount u32
	pStripeInfos    &RenderPassStripeInfoARM
}

// RenderPassStripeSubmitInfoARM extends VkCommandBufferSubmitInfo
pub type RenderPassStripeSubmitInfoARM = C.VkRenderPassStripeSubmitInfoARM

@[typedef]
pub struct C.VkRenderPassStripeSubmitInfoARM {
pub mut:
	sType                    StructureType = StructureType.render_pass_stripe_submit_info_arm
	pNext                    voidptr       = unsafe { nil }
	stripeSemaphoreInfoCount u32
	pStripeSemaphoreInfos    &SemaphoreSubmitInfo
}

pub const qcom_fragment_density_map_offset_spec_version = 3
pub const qcom_fragment_density_map_offset_extension_name = c'VK_QCOM_fragment_density_map_offset'
// PhysicalDeviceFragmentDensityMapOffsetFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceFragmentDensityMapOffsetFeaturesEXT = C.VkPhysicalDeviceFragmentDensityMapOffsetFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceFragmentDensityMapOffsetFeaturesEXT {
pub mut:
	sType                    StructureType = StructureType.physical_device_fragment_density_map_offset_features_ext
	pNext                    voidptr       = unsafe { nil }
	fragmentDensityMapOffset Bool32
}

pub type PhysicalDeviceFragmentDensityMapOffsetFeaturesQCOM = C.VkPhysicalDeviceFragmentDensityMapOffsetFeaturesEXT

// PhysicalDeviceFragmentDensityMapOffsetPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceFragmentDensityMapOffsetPropertiesEXT = C.VkPhysicalDeviceFragmentDensityMapOffsetPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceFragmentDensityMapOffsetPropertiesEXT {
pub mut:
	sType                            StructureType = StructureType.physical_device_fragment_density_map_offset_properties_ext
	pNext                            voidptr       = unsafe { nil }
	fragmentDensityOffsetGranularity Extent2D
}

pub type PhysicalDeviceFragmentDensityMapOffsetPropertiesQCOM = C.VkPhysicalDeviceFragmentDensityMapOffsetPropertiesEXT

// RenderPassFragmentDensityMapOffsetEndInfoEXT extends VkSubpassEndInfo,VkRenderingEndInfoKHR
pub type RenderPassFragmentDensityMapOffsetEndInfoEXT = C.VkRenderPassFragmentDensityMapOffsetEndInfoEXT

@[typedef]
pub struct C.VkRenderPassFragmentDensityMapOffsetEndInfoEXT {
pub mut:
	sType                      StructureType = StructureType.render_pass_fragment_density_map_offset_end_info_ext
	pNext                      voidptr       = unsafe { nil }
	fragmentDensityOffsetCount u32
	pFragmentDensityOffsets    &Offset2D
}

pub type SubpassFragmentDensityMapOffsetEndInfoQCOM = C.VkRenderPassFragmentDensityMapOffsetEndInfoEXT

pub const nv_copy_memory_indirect_spec_version = 1
pub const nv_copy_memory_indirect_extension_name = c'VK_NV_copy_memory_indirect'

pub type CopyMemoryIndirectCommandNV = C.VkCopyMemoryIndirectCommandKHR

pub type CopyMemoryToImageIndirectCommandNV = C.VkCopyMemoryToImageIndirectCommandKHR

// PhysicalDeviceCopyMemoryIndirectFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCopyMemoryIndirectFeaturesNV = C.VkPhysicalDeviceCopyMemoryIndirectFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceCopyMemoryIndirectFeaturesNV {
pub mut:
	sType        StructureType = StructureType.physical_device_copy_memory_indirect_features_nv
	pNext        voidptr       = unsafe { nil }
	indirectCopy Bool32
}

pub type PhysicalDeviceCopyMemoryIndirectPropertiesNV = C.VkPhysicalDeviceCopyMemoryIndirectPropertiesKHR

@[keep_args_alive]
fn C.vkCmdCopyMemoryIndirectNV(command_buffer CommandBuffer, copy_buffer_address DeviceAddress, copy_count u32, stride u32)

pub type PFN_vkCmdCopyMemoryIndirectNV = fn (command_buffer CommandBuffer, copy_buffer_address DeviceAddress, copy_count u32, stride u32)

@[inline]
pub fn cmd_copy_memory_indirect_nv(command_buffer CommandBuffer,
	copy_buffer_address DeviceAddress,
	copy_count u32,
	stride u32) {
	C.vkCmdCopyMemoryIndirectNV(command_buffer, copy_buffer_address, copy_count, stride)
}

@[keep_args_alive]
fn C.vkCmdCopyMemoryToImageIndirectNV(command_buffer CommandBuffer, copy_buffer_address DeviceAddress, copy_count u32, stride u32, dst_image Image, dst_image_layout ImageLayout, p_image_subresources &ImageSubresourceLayers)

pub type PFN_vkCmdCopyMemoryToImageIndirectNV = fn (command_buffer CommandBuffer, copy_buffer_address DeviceAddress, copy_count u32, stride u32, dst_image Image, dst_image_layout ImageLayout, p_image_subresources &ImageSubresourceLayers)

@[inline]
pub fn cmd_copy_memory_to_image_indirect_nv(command_buffer CommandBuffer,
	copy_buffer_address DeviceAddress,
	copy_count u32,
	stride u32,
	dst_image Image,
	dst_image_layout ImageLayout,
	p_image_subresources &ImageSubresourceLayers) {
	C.vkCmdCopyMemoryToImageIndirectNV(command_buffer, copy_buffer_address, copy_count,
		stride, dst_image, dst_image_layout, p_image_subresources)
}

pub const nv_memory_decompression_spec_version = 1
pub const nv_memory_decompression_extension_name = c'VK_NV_memory_decompression'

// Flag bits for MemoryDecompressionMethodFlagBitsEXT
pub type MemoryDecompressionMethodFlagBitsEXT = u64

pub const memory_decompression_method_gdeflate_1_0_bit_ext = u64(0x00000001)
pub const memory_decompression_method_gdeflate_1_0_bit_nv = memory_decompression_method_gdeflate_1_0_bit_ext

pub type MemoryDecompressionMethodFlagBitsNV = u64

pub type MemoryDecompressionMethodFlagsEXT = u64
pub type MemoryDecompressionMethodFlagsNV = u64
pub type DecompressMemoryRegionNV = C.VkDecompressMemoryRegionNV

@[typedef]
pub struct C.VkDecompressMemoryRegionNV {
pub mut:
	srcAddress          DeviceAddress
	dstAddress          DeviceAddress
	compressedSize      DeviceSize
	decompressedSize    DeviceSize
	decompressionMethod MemoryDecompressionMethodFlagsNV
}

// PhysicalDeviceMemoryDecompressionFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMemoryDecompressionFeaturesEXT = C.VkPhysicalDeviceMemoryDecompressionFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMemoryDecompressionFeaturesEXT {
pub mut:
	sType               StructureType = StructureType.physical_device_memory_decompression_features_ext
	pNext               voidptr       = unsafe { nil }
	memoryDecompression Bool32
}

pub type PhysicalDeviceMemoryDecompressionFeaturesNV = C.VkPhysicalDeviceMemoryDecompressionFeaturesEXT

// PhysicalDeviceMemoryDecompressionPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMemoryDecompressionPropertiesEXT = C.VkPhysicalDeviceMemoryDecompressionPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMemoryDecompressionPropertiesEXT {
pub mut:
	sType                         StructureType = StructureType.physical_device_memory_decompression_properties_ext
	pNext                         voidptr       = unsafe { nil }
	decompressionMethods          MemoryDecompressionMethodFlagsEXT
	maxDecompressionIndirectCount u64
}

pub type PhysicalDeviceMemoryDecompressionPropertiesNV = C.VkPhysicalDeviceMemoryDecompressionPropertiesEXT

@[keep_args_alive]
fn C.vkCmdDecompressMemoryNV(command_buffer CommandBuffer, decompress_region_count u32, p_decompress_memory_regions &DecompressMemoryRegionNV)

pub type PFN_vkCmdDecompressMemoryNV = fn (command_buffer CommandBuffer, decompress_region_count u32, p_decompress_memory_regions &DecompressMemoryRegionNV)

@[inline]
pub fn cmd_decompress_memory_nv(command_buffer CommandBuffer,
	decompress_region_count u32,
	p_decompress_memory_regions &DecompressMemoryRegionNV) {
	C.vkCmdDecompressMemoryNV(command_buffer, decompress_region_count, p_decompress_memory_regions)
}

@[keep_args_alive]
fn C.vkCmdDecompressMemoryIndirectCountNV(command_buffer CommandBuffer, indirect_commands_address DeviceAddress, indirect_commands_count_address DeviceAddress, stride u32)

pub type PFN_vkCmdDecompressMemoryIndirectCountNV = fn (command_buffer CommandBuffer, indirect_commands_address DeviceAddress, indirect_commands_count_address DeviceAddress, stride u32)

@[inline]
pub fn cmd_decompress_memory_indirect_count_nv(command_buffer CommandBuffer,
	indirect_commands_address DeviceAddress,
	indirect_commands_count_address DeviceAddress,
	stride u32) {
	C.vkCmdDecompressMemoryIndirectCountNV(command_buffer, indirect_commands_address,
		indirect_commands_count_address, stride)
}

pub const nv_device_generated_commands_compute_spec_version = 2
pub const nv_device_generated_commands_compute_extension_name = c'VK_NV_device_generated_commands_compute'
// PhysicalDeviceDeviceGeneratedCommandsComputeFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDeviceGeneratedCommandsComputeFeaturesNV = C.VkPhysicalDeviceDeviceGeneratedCommandsComputeFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceDeviceGeneratedCommandsComputeFeaturesNV {
pub mut:
	sType                               StructureType = StructureType.physical_device_device_generated_commands_compute_features_nv
	pNext                               voidptr       = unsafe { nil }
	deviceGeneratedCompute              Bool32
	deviceGeneratedComputePipelines     Bool32
	deviceGeneratedComputeCaptureReplay Bool32
}

// ComputePipelineIndirectBufferInfoNV extends VkComputePipelineCreateInfo
pub type ComputePipelineIndirectBufferInfoNV = C.VkComputePipelineIndirectBufferInfoNV

@[typedef]
pub struct C.VkComputePipelineIndirectBufferInfoNV {
pub mut:
	sType                              StructureType = StructureType.compute_pipeline_indirect_buffer_info_nv
	pNext                              voidptr       = unsafe { nil }
	deviceAddress                      DeviceAddress
	size                               DeviceSize
	pipelineDeviceAddressCaptureReplay DeviceAddress
}

pub type PipelineIndirectDeviceAddressInfoNV = C.VkPipelineIndirectDeviceAddressInfoNV

@[typedef]
pub struct C.VkPipelineIndirectDeviceAddressInfoNV {
pub mut:
	sType             StructureType = StructureType.pipeline_indirect_device_address_info_nv
	pNext             voidptr       = unsafe { nil }
	pipelineBindPoint PipelineBindPoint
	pipeline          Pipeline
}

pub type BindPipelineIndirectCommandNV = C.VkBindPipelineIndirectCommandNV

@[typedef]
pub struct C.VkBindPipelineIndirectCommandNV {
pub mut:
	pipelineAddress DeviceAddress
}

@[keep_args_alive]
fn C.vkGetPipelineIndirectMemoryRequirementsNV(device Device, p_create_info &ComputePipelineCreateInfo, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetPipelineIndirectMemoryRequirementsNV = fn (device Device, p_create_info &ComputePipelineCreateInfo, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_pipeline_indirect_memory_requirements_nv(device Device,
	p_create_info &ComputePipelineCreateInfo,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetPipelineIndirectMemoryRequirementsNV(device, p_create_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkCmdUpdatePipelineIndirectBufferNV(command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, pipeline Pipeline)

pub type PFN_vkCmdUpdatePipelineIndirectBufferNV = fn (command_buffer CommandBuffer, pipeline_bind_point PipelineBindPoint, pipeline Pipeline)

@[inline]
pub fn cmd_update_pipeline_indirect_buffer_nv(command_buffer CommandBuffer,
	pipeline_bind_point PipelineBindPoint,
	pipeline Pipeline) {
	C.vkCmdUpdatePipelineIndirectBufferNV(command_buffer, pipeline_bind_point, pipeline)
}

@[keep_args_alive]
fn C.vkGetPipelineIndirectDeviceAddressNV(device Device, p_info &PipelineIndirectDeviceAddressInfoNV) DeviceAddress

pub type PFN_vkGetPipelineIndirectDeviceAddressNV = fn (device Device, p_info &PipelineIndirectDeviceAddressInfoNV) DeviceAddress

@[inline]
pub fn get_pipeline_indirect_device_address_nv(device Device,
	p_info &PipelineIndirectDeviceAddressInfoNV) DeviceAddress {
	return C.vkGetPipelineIndirectDeviceAddressNV(device, p_info)
}

pub const nv_ray_tracing_linear_swept_spheres_spec_version = 1
pub const nv_ray_tracing_linear_swept_spheres_extension_name = c'VK_NV_ray_tracing_linear_swept_spheres'

pub enum RayTracingLssIndexingModeNV as u32 {
	list        = 0
	successive  = 1
	max_enum_nv = max_int
}

pub enum RayTracingLssPrimitiveEndCapsModeNV as u32 {
	none        = 0
	chained     = 1
	max_enum_nv = max_int
}
// PhysicalDeviceRayTracingLinearSweptSpheresFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRayTracingLinearSweptSpheresFeaturesNV = C.VkPhysicalDeviceRayTracingLinearSweptSpheresFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceRayTracingLinearSweptSpheresFeaturesNV {
pub mut:
	sType              StructureType = StructureType.physical_device_ray_tracing_linear_swept_spheres_features_nv
	pNext              voidptr       = unsafe { nil }
	spheres            Bool32
	linearSweptSpheres Bool32
}

// AccelerationStructureGeometryLinearSweptSpheresDataNV extends VkAccelerationStructureGeometryKHR
pub type AccelerationStructureGeometryLinearSweptSpheresDataNV = C.VkAccelerationStructureGeometryLinearSweptSpheresDataNV

@[typedef]
pub struct C.VkAccelerationStructureGeometryLinearSweptSpheresDataNV {
pub mut:
	sType        StructureType = StructureType.acceleration_structure_geometry_linear_swept_spheres_data_nv
	pNext        voidptr       = unsafe { nil }
	vertexFormat Format
	vertexData   DeviceOrHostAddressConstKHR
	vertexStride DeviceSize
	radiusFormat Format
	radiusData   DeviceOrHostAddressConstKHR
	radiusStride DeviceSize
	indexType    IndexType
	indexData    DeviceOrHostAddressConstKHR
	indexStride  DeviceSize
	indexingMode RayTracingLssIndexingModeNV
	endCapsMode  RayTracingLssPrimitiveEndCapsModeNV
}

// AccelerationStructureGeometrySpheresDataNV extends VkAccelerationStructureGeometryKHR
pub type AccelerationStructureGeometrySpheresDataNV = C.VkAccelerationStructureGeometrySpheresDataNV

@[typedef]
pub struct C.VkAccelerationStructureGeometrySpheresDataNV {
pub mut:
	sType        StructureType = StructureType.acceleration_structure_geometry_spheres_data_nv
	pNext        voidptr       = unsafe { nil }
	vertexFormat Format
	vertexData   DeviceOrHostAddressConstKHR
	vertexStride DeviceSize
	radiusFormat Format
	radiusData   DeviceOrHostAddressConstKHR
	radiusStride DeviceSize
	indexType    IndexType
	indexData    DeviceOrHostAddressConstKHR
	indexStride  DeviceSize
}

pub const nv_linear_color_attachment_spec_version = 1
pub const nv_linear_color_attachment_extension_name = c'VK_NV_linear_color_attachment'
// PhysicalDeviceLinearColorAttachmentFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceLinearColorAttachmentFeaturesNV = C.VkPhysicalDeviceLinearColorAttachmentFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceLinearColorAttachmentFeaturesNV {
pub mut:
	sType                 StructureType = StructureType.physical_device_linear_color_attachment_features_nv
	pNext                 voidptr       = unsafe { nil }
	linearColorAttachment Bool32
}

pub const google_surfaceless_query_spec_version = 2
pub const google_surfaceless_query_extension_name = c'VK_GOOGE_surfaceless_query'

pub const ext_image_compression_control_swapchain_spec_version = 1
pub const ext_image_compression_control_swapchain_extension_name = c'VK_EXT_image_compression_control_swapchain'
// PhysicalDeviceImageCompressionControlSwapchainFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceImageCompressionControlSwapchainFeaturesEXT = C.VkPhysicalDeviceImageCompressionControlSwapchainFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceImageCompressionControlSwapchainFeaturesEXT {
pub mut:
	sType                            StructureType = StructureType.physical_device_image_compression_control_swapchain_features_ext
	pNext                            voidptr       = unsafe { nil }
	imageCompressionControlSwapchain Bool32
}

pub const qcom_image_processing_spec_version = 1
pub const qcom_image_processing_extension_name = c'VK_QCOM_image_processing'
// ImageViewSampleWeightCreateInfoQCOM extends VkImageViewCreateInfo
pub type ImageViewSampleWeightCreateInfoQCOM = C.VkImageViewSampleWeightCreateInfoQCOM

@[typedef]
pub struct C.VkImageViewSampleWeightCreateInfoQCOM {
pub mut:
	sType        StructureType = StructureType.image_view_sample_weight_create_info_qcom
	pNext        voidptr       = unsafe { nil }
	filterCenter Offset2D
	filterSize   Extent2D
	numPhases    u32
}

// PhysicalDeviceImageProcessingFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceImageProcessingFeaturesQCOM = C.VkPhysicalDeviceImageProcessingFeaturesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceImageProcessingFeaturesQCOM {
pub mut:
	sType                 StructureType = StructureType.physical_device_image_processing_features_qcom
	pNext                 voidptr       = unsafe { nil }
	textureSampleWeighted Bool32
	textureBoxFilter      Bool32
	textureBlockMatch     Bool32
}

// PhysicalDeviceImageProcessingPropertiesQCOM extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceImageProcessingPropertiesQCOM = C.VkPhysicalDeviceImageProcessingPropertiesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceImageProcessingPropertiesQCOM {
pub mut:
	sType                    StructureType = StructureType.physical_device_image_processing_properties_qcom
	pNext                    voidptr       = unsafe { nil }
	maxWeightFilterPhases    u32
	maxWeightFilterDimension Extent2D
	maxBlockMatchRegion      Extent2D
	maxBoxFilterBlockSize    Extent2D
}

pub const ext_nested_command_buffer_spec_version = 1
pub const ext_nested_command_buffer_extension_name = c'VK_EXT_nested_command_buffer'
// PhysicalDeviceNestedCommandBufferFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceNestedCommandBufferFeaturesEXT = C.VkPhysicalDeviceNestedCommandBufferFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceNestedCommandBufferFeaturesEXT {
pub mut:
	sType                              StructureType = StructureType.physical_device_nested_command_buffer_features_ext
	pNext                              voidptr       = unsafe { nil }
	nestedCommandBuffer                Bool32
	nestedCommandBufferRendering       Bool32
	nestedCommandBufferSimultaneousUse Bool32
}

// PhysicalDeviceNestedCommandBufferPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceNestedCommandBufferPropertiesEXT = C.VkPhysicalDeviceNestedCommandBufferPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceNestedCommandBufferPropertiesEXT {
pub mut:
	sType                        StructureType = StructureType.physical_device_nested_command_buffer_properties_ext
	pNext                        voidptr       = unsafe { nil }
	maxCommandBufferNestingLevel u32
}

pub const ext_external_memory_acquire_unmodified_spec_version = 1
pub const ext_external_memory_acquire_unmodified_extension_name = c'VK_EXT_external_memory_acquire_unmodified'
// ExternalMemoryAcquireUnmodifiedEXT extends VkBufferMemoryBarrier,VkBufferMemoryBarrier2,VkImageMemoryBarrier,VkImageMemoryBarrier2
pub type ExternalMemoryAcquireUnmodifiedEXT = C.VkExternalMemoryAcquireUnmodifiedEXT

@[typedef]
pub struct C.VkExternalMemoryAcquireUnmodifiedEXT {
pub mut:
	sType                   StructureType = StructureType.external_memory_acquire_unmodified_ext
	pNext                   voidptr       = unsafe { nil }
	acquireUnmodifiedMemory Bool32
}

pub const ext_extended_dynamic_state_3_spec_version = 2
pub const ext_extended_dynamic_state_3_extension_name = c'VK_EXT_extended_dynamic_state3'
// PhysicalDeviceExtendedDynamicState3FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceExtendedDynamicState3FeaturesEXT = C.VkPhysicalDeviceExtendedDynamicState3FeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceExtendedDynamicState3FeaturesEXT {
pub mut:
	sType                                                 StructureType = StructureType.physical_device_extended_dynamic_state3_features_ext
	pNext                                                 voidptr       = unsafe { nil }
	extendedDynamicState3TessellationDomainOrigin         Bool32
	extendedDynamicState3DepthClampEnable                 Bool32
	extendedDynamicState3PolygonMode                      Bool32
	extendedDynamicState3RasterizationSamples             Bool32
	extendedDynamicState3SampleMask                       Bool32
	extendedDynamicState3AlphaToCoverageEnable            Bool32
	extendedDynamicState3AlphaToOneEnable                 Bool32
	extendedDynamicState3LogicOpEnable                    Bool32
	extendedDynamicState3ColorBlendEnable                 Bool32
	extendedDynamicState3ColorBlendEquation               Bool32
	extendedDynamicState3ColorWriteMask                   Bool32
	extendedDynamicState3RasterizationStream              Bool32
	extendedDynamicState3ConservativeRasterizationMode    Bool32
	extendedDynamicState3ExtraPrimitiveOverestimationSize Bool32
	extendedDynamicState3DepthClipEnable                  Bool32
	extendedDynamicState3SampleLocationsEnable            Bool32
	extendedDynamicState3ColorBlendAdvanced               Bool32
	extendedDynamicState3ProvokingVertexMode              Bool32
	extendedDynamicState3LineRasterizationMode            Bool32
	extendedDynamicState3LineStippleEnable                Bool32
	extendedDynamicState3DepthClipNegativeOneToOne        Bool32
	extendedDynamicState3ViewportWScalingEnable           Bool32
	extendedDynamicState3ViewportSwizzle                  Bool32
	extendedDynamicState3CoverageToColorEnable            Bool32
	extendedDynamicState3CoverageToColorLocation          Bool32
	extendedDynamicState3CoverageModulationMode           Bool32
	extendedDynamicState3CoverageModulationTableEnable    Bool32
	extendedDynamicState3CoverageModulationTable          Bool32
	extendedDynamicState3CoverageReductionMode            Bool32
	extendedDynamicState3RepresentativeFragmentTestEnable Bool32
	extendedDynamicState3ShadingRateImageEnable           Bool32
}

// PhysicalDeviceExtendedDynamicState3PropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceExtendedDynamicState3PropertiesEXT = C.VkPhysicalDeviceExtendedDynamicState3PropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceExtendedDynamicState3PropertiesEXT {
pub mut:
	sType                                StructureType = StructureType.physical_device_extended_dynamic_state3_properties_ext
	pNext                                voidptr       = unsafe { nil }
	dynamicPrimitiveTopologyUnrestricted Bool32
}

pub type ColorBlendEquationEXT = C.VkColorBlendEquationEXT

@[typedef]
pub struct C.VkColorBlendEquationEXT {
pub mut:
	srcColorBlendFactor BlendFactor
	dstColorBlendFactor BlendFactor
	colorBlendOp        BlendOp
	srcAlphaBlendFactor BlendFactor
	dstAlphaBlendFactor BlendFactor
	alphaBlendOp        BlendOp
}

pub type ColorBlendAdvancedEXT = C.VkColorBlendAdvancedEXT

@[typedef]
pub struct C.VkColorBlendAdvancedEXT {
pub mut:
	advancedBlendOp  BlendOp
	srcPremultiplied Bool32
	dstPremultiplied Bool32
	blendOverlap     BlendOverlapEXT
	clampResults     Bool32
}

@[keep_args_alive]
fn C.vkCmdSetDepthClampEnableEXT(command_buffer CommandBuffer, depth_clamp_enable Bool32)

pub type PFN_vkCmdSetDepthClampEnableEXT = fn (command_buffer CommandBuffer, depth_clamp_enable Bool32)

@[inline]
pub fn cmd_set_depth_clamp_enable_ext(command_buffer CommandBuffer,
	depth_clamp_enable Bool32) {
	C.vkCmdSetDepthClampEnableEXT(command_buffer, depth_clamp_enable)
}

@[keep_args_alive]
fn C.vkCmdSetPolygonModeEXT(command_buffer CommandBuffer, polygon_mode PolygonMode)

pub type PFN_vkCmdSetPolygonModeEXT = fn (command_buffer CommandBuffer, polygon_mode PolygonMode)

@[inline]
pub fn cmd_set_polygon_mode_ext(command_buffer CommandBuffer,
	polygon_mode PolygonMode) {
	C.vkCmdSetPolygonModeEXT(command_buffer, polygon_mode)
}

@[keep_args_alive]
fn C.vkCmdSetRasterizationSamplesEXT(command_buffer CommandBuffer, rasterization_samples SampleCountFlagBits)

pub type PFN_vkCmdSetRasterizationSamplesEXT = fn (command_buffer CommandBuffer, rasterization_samples SampleCountFlagBits)

@[inline]
pub fn cmd_set_rasterization_samples_ext(command_buffer CommandBuffer,
	rasterization_samples SampleCountFlagBits) {
	C.vkCmdSetRasterizationSamplesEXT(command_buffer, rasterization_samples)
}

@[keep_args_alive]
fn C.vkCmdSetSampleMaskEXT(command_buffer CommandBuffer, samples SampleCountFlagBits, p_sample_mask &SampleMask)

pub type PFN_vkCmdSetSampleMaskEXT = fn (command_buffer CommandBuffer, samples SampleCountFlagBits, p_sample_mask &SampleMask)

@[inline]
pub fn cmd_set_sample_mask_ext(command_buffer CommandBuffer,
	samples SampleCountFlagBits,
	p_sample_mask &SampleMask) {
	C.vkCmdSetSampleMaskEXT(command_buffer, samples, p_sample_mask)
}

@[keep_args_alive]
fn C.vkCmdSetAlphaToCoverageEnableEXT(command_buffer CommandBuffer, alpha_to_coverage_enable Bool32)

pub type PFN_vkCmdSetAlphaToCoverageEnableEXT = fn (command_buffer CommandBuffer, alpha_to_coverage_enable Bool32)

@[inline]
pub fn cmd_set_alpha_to_coverage_enable_ext(command_buffer CommandBuffer,
	alpha_to_coverage_enable Bool32) {
	C.vkCmdSetAlphaToCoverageEnableEXT(command_buffer, alpha_to_coverage_enable)
}

@[keep_args_alive]
fn C.vkCmdSetAlphaToOneEnableEXT(command_buffer CommandBuffer, alpha_to_one_enable Bool32)

pub type PFN_vkCmdSetAlphaToOneEnableEXT = fn (command_buffer CommandBuffer, alpha_to_one_enable Bool32)

@[inline]
pub fn cmd_set_alpha_to_one_enable_ext(command_buffer CommandBuffer,
	alpha_to_one_enable Bool32) {
	C.vkCmdSetAlphaToOneEnableEXT(command_buffer, alpha_to_one_enable)
}

@[keep_args_alive]
fn C.vkCmdSetLogicOpEnableEXT(command_buffer CommandBuffer, logic_op_enable Bool32)

pub type PFN_vkCmdSetLogicOpEnableEXT = fn (command_buffer CommandBuffer, logic_op_enable Bool32)

@[inline]
pub fn cmd_set_logic_op_enable_ext(command_buffer CommandBuffer,
	logic_op_enable Bool32) {
	C.vkCmdSetLogicOpEnableEXT(command_buffer, logic_op_enable)
}

@[keep_args_alive]
fn C.vkCmdSetColorBlendEnableEXT(command_buffer CommandBuffer, first_attachment u32, attachment_count u32, p_color_blend_enables &Bool32)

pub type PFN_vkCmdSetColorBlendEnableEXT = fn (command_buffer CommandBuffer, first_attachment u32, attachment_count u32, p_color_blend_enables &Bool32)

@[inline]
pub fn cmd_set_color_blend_enable_ext(command_buffer CommandBuffer,
	first_attachment u32,
	attachment_count u32,
	p_color_blend_enables &Bool32) {
	C.vkCmdSetColorBlendEnableEXT(command_buffer, first_attachment, attachment_count,
		p_color_blend_enables)
}

@[keep_args_alive]
fn C.vkCmdSetColorBlendEquationEXT(command_buffer CommandBuffer, first_attachment u32, attachment_count u32, p_color_blend_equations &ColorBlendEquationEXT)

pub type PFN_vkCmdSetColorBlendEquationEXT = fn (command_buffer CommandBuffer, first_attachment u32, attachment_count u32, p_color_blend_equations &ColorBlendEquationEXT)

@[inline]
pub fn cmd_set_color_blend_equation_ext(command_buffer CommandBuffer,
	first_attachment u32,
	attachment_count u32,
	p_color_blend_equations &ColorBlendEquationEXT) {
	C.vkCmdSetColorBlendEquationEXT(command_buffer, first_attachment, attachment_count,
		p_color_blend_equations)
}

@[keep_args_alive]
fn C.vkCmdSetColorWriteMaskEXT(command_buffer CommandBuffer, first_attachment u32, attachment_count u32, p_color_write_masks &ColorComponentFlags)

pub type PFN_vkCmdSetColorWriteMaskEXT = fn (command_buffer CommandBuffer, first_attachment u32, attachment_count u32, p_color_write_masks &ColorComponentFlags)

@[inline]
pub fn cmd_set_color_write_mask_ext(command_buffer CommandBuffer,
	first_attachment u32,
	attachment_count u32,
	p_color_write_masks &ColorComponentFlags) {
	C.vkCmdSetColorWriteMaskEXT(command_buffer, first_attachment, attachment_count, p_color_write_masks)
}

@[keep_args_alive]
fn C.vkCmdSetTessellationDomainOriginEXT(command_buffer CommandBuffer, domain_origin TessellationDomainOrigin)

pub type PFN_vkCmdSetTessellationDomainOriginEXT = fn (command_buffer CommandBuffer, domain_origin TessellationDomainOrigin)

@[inline]
pub fn cmd_set_tessellation_domain_origin_ext(command_buffer CommandBuffer,
	domain_origin TessellationDomainOrigin) {
	C.vkCmdSetTessellationDomainOriginEXT(command_buffer, domain_origin)
}

@[keep_args_alive]
fn C.vkCmdSetRasterizationStreamEXT(command_buffer CommandBuffer, rasterization_stream u32)

pub type PFN_vkCmdSetRasterizationStreamEXT = fn (command_buffer CommandBuffer, rasterization_stream u32)

@[inline]
pub fn cmd_set_rasterization_stream_ext(command_buffer CommandBuffer,
	rasterization_stream u32) {
	C.vkCmdSetRasterizationStreamEXT(command_buffer, rasterization_stream)
}

@[keep_args_alive]
fn C.vkCmdSetConservativeRasterizationModeEXT(command_buffer CommandBuffer, conservative_rasterization_mode ConservativeRasterizationModeEXT)

pub type PFN_vkCmdSetConservativeRasterizationModeEXT = fn (command_buffer CommandBuffer, conservative_rasterization_mode ConservativeRasterizationModeEXT)

@[inline]
pub fn cmd_set_conservative_rasterization_mode_ext(command_buffer CommandBuffer,
	conservative_rasterization_mode ConservativeRasterizationModeEXT) {
	C.vkCmdSetConservativeRasterizationModeEXT(command_buffer, conservative_rasterization_mode)
}

@[keep_args_alive]
fn C.vkCmdSetExtraPrimitiveOverestimationSizeEXT(command_buffer CommandBuffer, extra_primitive_overestimation_size f32)

pub type PFN_vkCmdSetExtraPrimitiveOverestimationSizeEXT = fn (command_buffer CommandBuffer, extra_primitive_overestimation_size f32)

@[inline]
pub fn cmd_set_extra_primitive_overestimation_size_ext(command_buffer CommandBuffer,
	extra_primitive_overestimation_size f32) {
	C.vkCmdSetExtraPrimitiveOverestimationSizeEXT(command_buffer, extra_primitive_overestimation_size)
}

@[keep_args_alive]
fn C.vkCmdSetDepthClipEnableEXT(command_buffer CommandBuffer, depth_clip_enable Bool32)

pub type PFN_vkCmdSetDepthClipEnableEXT = fn (command_buffer CommandBuffer, depth_clip_enable Bool32)

@[inline]
pub fn cmd_set_depth_clip_enable_ext(command_buffer CommandBuffer,
	depth_clip_enable Bool32) {
	C.vkCmdSetDepthClipEnableEXT(command_buffer, depth_clip_enable)
}

@[keep_args_alive]
fn C.vkCmdSetSampleLocationsEnableEXT(command_buffer CommandBuffer, sample_locations_enable Bool32)

pub type PFN_vkCmdSetSampleLocationsEnableEXT = fn (command_buffer CommandBuffer, sample_locations_enable Bool32)

@[inline]
pub fn cmd_set_sample_locations_enable_ext(command_buffer CommandBuffer,
	sample_locations_enable Bool32) {
	C.vkCmdSetSampleLocationsEnableEXT(command_buffer, sample_locations_enable)
}

@[keep_args_alive]
fn C.vkCmdSetColorBlendAdvancedEXT(command_buffer CommandBuffer, first_attachment u32, attachment_count u32, p_color_blend_advanced &ColorBlendAdvancedEXT)

pub type PFN_vkCmdSetColorBlendAdvancedEXT = fn (command_buffer CommandBuffer, first_attachment u32, attachment_count u32, p_color_blend_advanced &ColorBlendAdvancedEXT)

@[inline]
pub fn cmd_set_color_blend_advanced_ext(command_buffer CommandBuffer,
	first_attachment u32,
	attachment_count u32,
	p_color_blend_advanced &ColorBlendAdvancedEXT) {
	C.vkCmdSetColorBlendAdvancedEXT(command_buffer, first_attachment, attachment_count,
		p_color_blend_advanced)
}

@[keep_args_alive]
fn C.vkCmdSetProvokingVertexModeEXT(command_buffer CommandBuffer, provoking_vertex_mode ProvokingVertexModeEXT)

pub type PFN_vkCmdSetProvokingVertexModeEXT = fn (command_buffer CommandBuffer, provoking_vertex_mode ProvokingVertexModeEXT)

@[inline]
pub fn cmd_set_provoking_vertex_mode_ext(command_buffer CommandBuffer,
	provoking_vertex_mode ProvokingVertexModeEXT) {
	C.vkCmdSetProvokingVertexModeEXT(command_buffer, provoking_vertex_mode)
}

@[keep_args_alive]
fn C.vkCmdSetLineRasterizationModeEXT(command_buffer CommandBuffer, line_rasterization_mode LineRasterizationModeEXT)

pub type PFN_vkCmdSetLineRasterizationModeEXT = fn (command_buffer CommandBuffer, line_rasterization_mode LineRasterizationModeEXT)

@[inline]
pub fn cmd_set_line_rasterization_mode_ext(command_buffer CommandBuffer,
	line_rasterization_mode LineRasterizationModeEXT) {
	C.vkCmdSetLineRasterizationModeEXT(command_buffer, line_rasterization_mode)
}

@[keep_args_alive]
fn C.vkCmdSetLineStippleEnableEXT(command_buffer CommandBuffer, stippled_line_enable Bool32)

pub type PFN_vkCmdSetLineStippleEnableEXT = fn (command_buffer CommandBuffer, stippled_line_enable Bool32)

@[inline]
pub fn cmd_set_line_stipple_enable_ext(command_buffer CommandBuffer,
	stippled_line_enable Bool32) {
	C.vkCmdSetLineStippleEnableEXT(command_buffer, stippled_line_enable)
}

@[keep_args_alive]
fn C.vkCmdSetDepthClipNegativeOneToOneEXT(command_buffer CommandBuffer, negative_one_to_one Bool32)

pub type PFN_vkCmdSetDepthClipNegativeOneToOneEXT = fn (command_buffer CommandBuffer, negative_one_to_one Bool32)

@[inline]
pub fn cmd_set_depth_clip_negative_one_to_one_ext(command_buffer CommandBuffer,
	negative_one_to_one Bool32) {
	C.vkCmdSetDepthClipNegativeOneToOneEXT(command_buffer, negative_one_to_one)
}

@[keep_args_alive]
fn C.vkCmdSetViewportWScalingEnableNV(command_buffer CommandBuffer, viewport_w_scaling_enable Bool32)

pub type PFN_vkCmdSetViewportWScalingEnableNV = fn (command_buffer CommandBuffer, viewport_w_scaling_enable Bool32)

@[inline]
pub fn cmd_set_viewport_w_scaling_enable_nv(command_buffer CommandBuffer,
	viewport_w_scaling_enable Bool32) {
	C.vkCmdSetViewportWScalingEnableNV(command_buffer, viewport_w_scaling_enable)
}

@[keep_args_alive]
fn C.vkCmdSetViewportSwizzleNV(command_buffer CommandBuffer, first_viewport u32, viewport_count u32, p_viewport_swizzles &ViewportSwizzleNV)

pub type PFN_vkCmdSetViewportSwizzleNV = fn (command_buffer CommandBuffer, first_viewport u32, viewport_count u32, p_viewport_swizzles &ViewportSwizzleNV)

@[inline]
pub fn cmd_set_viewport_swizzle_nv(command_buffer CommandBuffer,
	first_viewport u32,
	viewport_count u32,
	p_viewport_swizzles &ViewportSwizzleNV) {
	C.vkCmdSetViewportSwizzleNV(command_buffer, first_viewport, viewport_count, p_viewport_swizzles)
}

@[keep_args_alive]
fn C.vkCmdSetCoverageToColorEnableNV(command_buffer CommandBuffer, coverage_to_color_enable Bool32)

pub type PFN_vkCmdSetCoverageToColorEnableNV = fn (command_buffer CommandBuffer, coverage_to_color_enable Bool32)

@[inline]
pub fn cmd_set_coverage_to_color_enable_nv(command_buffer CommandBuffer,
	coverage_to_color_enable Bool32) {
	C.vkCmdSetCoverageToColorEnableNV(command_buffer, coverage_to_color_enable)
}

@[keep_args_alive]
fn C.vkCmdSetCoverageToColorLocationNV(command_buffer CommandBuffer, coverage_to_color_location u32)

pub type PFN_vkCmdSetCoverageToColorLocationNV = fn (command_buffer CommandBuffer, coverage_to_color_location u32)

@[inline]
pub fn cmd_set_coverage_to_color_location_nv(command_buffer CommandBuffer,
	coverage_to_color_location u32) {
	C.vkCmdSetCoverageToColorLocationNV(command_buffer, coverage_to_color_location)
}

@[keep_args_alive]
fn C.vkCmdSetCoverageModulationModeNV(command_buffer CommandBuffer, coverage_modulation_mode CoverageModulationModeNV)

pub type PFN_vkCmdSetCoverageModulationModeNV = fn (command_buffer CommandBuffer, coverage_modulation_mode CoverageModulationModeNV)

@[inline]
pub fn cmd_set_coverage_modulation_mode_nv(command_buffer CommandBuffer,
	coverage_modulation_mode CoverageModulationModeNV) {
	C.vkCmdSetCoverageModulationModeNV(command_buffer, coverage_modulation_mode)
}

@[keep_args_alive]
fn C.vkCmdSetCoverageModulationTableEnableNV(command_buffer CommandBuffer, coverage_modulation_table_enable Bool32)

pub type PFN_vkCmdSetCoverageModulationTableEnableNV = fn (command_buffer CommandBuffer, coverage_modulation_table_enable Bool32)

@[inline]
pub fn cmd_set_coverage_modulation_table_enable_nv(command_buffer CommandBuffer,
	coverage_modulation_table_enable Bool32) {
	C.vkCmdSetCoverageModulationTableEnableNV(command_buffer, coverage_modulation_table_enable)
}

@[keep_args_alive]
fn C.vkCmdSetCoverageModulationTableNV(command_buffer CommandBuffer, coverage_modulation_table_count u32, p_coverage_modulation_table &f32)

pub type PFN_vkCmdSetCoverageModulationTableNV = fn (command_buffer CommandBuffer, coverage_modulation_table_count u32, p_coverage_modulation_table &f32)

@[inline]
pub fn cmd_set_coverage_modulation_table_nv(command_buffer CommandBuffer,
	coverage_modulation_table_count u32,
	p_coverage_modulation_table &f32) {
	C.vkCmdSetCoverageModulationTableNV(command_buffer, coverage_modulation_table_count,
		p_coverage_modulation_table)
}

@[keep_args_alive]
fn C.vkCmdSetShadingRateImageEnableNV(command_buffer CommandBuffer, shading_rate_image_enable Bool32)

pub type PFN_vkCmdSetShadingRateImageEnableNV = fn (command_buffer CommandBuffer, shading_rate_image_enable Bool32)

@[inline]
pub fn cmd_set_shading_rate_image_enable_nv(command_buffer CommandBuffer,
	shading_rate_image_enable Bool32) {
	C.vkCmdSetShadingRateImageEnableNV(command_buffer, shading_rate_image_enable)
}

@[keep_args_alive]
fn C.vkCmdSetRepresentativeFragmentTestEnableNV(command_buffer CommandBuffer, representative_fragment_test_enable Bool32)

pub type PFN_vkCmdSetRepresentativeFragmentTestEnableNV = fn (command_buffer CommandBuffer, representative_fragment_test_enable Bool32)

@[inline]
pub fn cmd_set_representative_fragment_test_enable_nv(command_buffer CommandBuffer,
	representative_fragment_test_enable Bool32) {
	C.vkCmdSetRepresentativeFragmentTestEnableNV(command_buffer, representative_fragment_test_enable)
}

@[keep_args_alive]
fn C.vkCmdSetCoverageReductionModeNV(command_buffer CommandBuffer, coverage_reduction_mode CoverageReductionModeNV)

pub type PFN_vkCmdSetCoverageReductionModeNV = fn (command_buffer CommandBuffer, coverage_reduction_mode CoverageReductionModeNV)

@[inline]
pub fn cmd_set_coverage_reduction_mode_nv(command_buffer CommandBuffer,
	coverage_reduction_mode CoverageReductionModeNV) {
	C.vkCmdSetCoverageReductionModeNV(command_buffer, coverage_reduction_mode)
}

pub const ext_subpass_merge_feedback_spec_version = 2
pub const ext_subpass_merge_feedback_extension_name = c'VK_EXT_subpass_merge_feedback'

pub enum SubpassMergeStatusEXT as u32 {
	merged                                   = 0
	disallowed                               = 1
	not_merged_side_effects                  = 2
	not_merged_samples_mismatch              = 3
	not_merged_views_mismatch                = 4
	not_merged_aliasing                      = 5
	not_merged_dependencies                  = 6
	not_merged_incompatible_input_attachment = 7
	not_merged_too_many_attachments          = 8
	not_merged_insufficient_storage          = 9
	not_merged_depth_stencil_count           = 10
	not_merged_resolve_attachment_reuse      = 11
	not_merged_single_subpass                = 12
	not_merged_unspecified                   = 13
	max_enum_ext                             = max_int
}
// PhysicalDeviceSubpassMergeFeedbackFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceSubpassMergeFeedbackFeaturesEXT = C.VkPhysicalDeviceSubpassMergeFeedbackFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceSubpassMergeFeedbackFeaturesEXT {
pub mut:
	sType                StructureType = StructureType.physical_device_subpass_merge_feedback_features_ext
	pNext                voidptr       = unsafe { nil }
	subpassMergeFeedback Bool32
}

// RenderPassCreationControlEXT extends VkRenderPassCreateInfo2,VkSubpassDescription2
pub type RenderPassCreationControlEXT = C.VkRenderPassCreationControlEXT

@[typedef]
pub struct C.VkRenderPassCreationControlEXT {
pub mut:
	sType           StructureType = StructureType.render_pass_creation_control_ext
	pNext           voidptr       = unsafe { nil }
	disallowMerging Bool32
}

pub type RenderPassCreationFeedbackInfoEXT = C.VkRenderPassCreationFeedbackInfoEXT

@[typedef]
pub struct C.VkRenderPassCreationFeedbackInfoEXT {
pub mut:
	postMergeSubpassCount u32
}

// RenderPassCreationFeedbackCreateInfoEXT extends VkRenderPassCreateInfo2
pub type RenderPassCreationFeedbackCreateInfoEXT = C.VkRenderPassCreationFeedbackCreateInfoEXT

@[typedef]
pub struct C.VkRenderPassCreationFeedbackCreateInfoEXT {
pub mut:
	sType               StructureType = StructureType.render_pass_creation_feedback_create_info_ext
	pNext               voidptr       = unsafe { nil }
	pRenderPassFeedback &RenderPassCreationFeedbackInfoEXT
}

pub type RenderPassSubpassFeedbackInfoEXT = C.VkRenderPassSubpassFeedbackInfoEXT

@[typedef]
pub struct C.VkRenderPassSubpassFeedbackInfoEXT {
pub mut:
	subpassMergeStatus SubpassMergeStatusEXT
	description        [max_description_size]char
	postMergeIndex     u32
}

// RenderPassSubpassFeedbackCreateInfoEXT extends VkSubpassDescription2
pub type RenderPassSubpassFeedbackCreateInfoEXT = C.VkRenderPassSubpassFeedbackCreateInfoEXT

@[typedef]
pub struct C.VkRenderPassSubpassFeedbackCreateInfoEXT {
pub mut:
	sType            StructureType = StructureType.render_pass_subpass_feedback_create_info_ext
	pNext            voidptr       = unsafe { nil }
	pSubpassFeedback &RenderPassSubpassFeedbackInfoEXT
}

pub const lunarg_direct_driver_loading_spec_version = 1
pub const lunarg_direct_driver_loading_extension_name = c'VK_NARG_direct_driver_loading'

pub enum DirectDriverLoadingModeLUNARG as u32 {
	exclusive       = 0
	inclusive       = 1
	max_enum_lunarg = max_int
}
pub type DirectDriverLoadingFlagsLUNARG = u32
pub type PFN_vkGetInstanceProcAddrLUNARG = fn (Instance, &char)

pub type DirectDriverLoadingInfoLUNARG = C.VkDirectDriverLoadingInfoLUNARG

@[typedef]
pub struct C.VkDirectDriverLoadingInfoLUNARG {
pub mut:
	sType                  StructureType = StructureType.direct_driver_loading_info_lunarg
	pNext                  voidptr       = unsafe { nil }
	flags                  DirectDriverLoadingFlagsLUNARG
	pfnGetInstanceProcAddr PFN_vkGetInstanceProcAddrLUNARG = unsafe { nil }
}

// DirectDriverLoadingListLUNARG extends VkInstanceCreateInfo
pub type DirectDriverLoadingListLUNARG = C.VkDirectDriverLoadingListLUNARG

@[typedef]
pub struct C.VkDirectDriverLoadingListLUNARG {
pub mut:
	sType       StructureType = StructureType.direct_driver_loading_list_lunarg
	pNext       voidptr       = unsafe { nil }
	mode        DirectDriverLoadingModeLUNARG
	driverCount u32
	pDrivers    &DirectDriverLoadingInfoLUNARG
}

// Pointer to VkTensorARM_T
pub type TensorARM = voidptr

// Pointer to VkTensorViewARM_T
pub type TensorViewARM = voidptr

pub const arm_tensors_spec_version = 1
pub const arm_tensors_extension_name = c'VK_ARM_tensors'

pub enum TensorTilingARM as u32 {
	optimal      = 0
	linear       = 1
	max_enum_arm = max_int
}
pub type TensorCreateFlagsARM = u64

// Flag bits for TensorCreateFlagBitsARM
pub type TensorCreateFlagBitsARM = u64

pub const tensor_create_mutable_format_bit_arm = u64(0x00000001)
pub const tensor_create_protected_bit_arm = u64(0x00000002)
pub const tensor_create_descriptor_buffer_capture_replay_bit_arm = u64(0x00000004)

pub type TensorViewCreateFlagsARM = u64

// Flag bits for TensorViewCreateFlagBitsARM
pub type TensorViewCreateFlagBitsARM = u64

pub const tensor_view_create_descriptor_buffer_capture_replay_bit_arm = u64(0x00000001)

pub type TensorUsageFlagsARM = u64

// Flag bits for TensorUsageFlagBitsARM
pub type TensorUsageFlagBitsARM = u64

pub const tensor_usage_shader_bit_arm = u64(0x00000002)
pub const tensor_usage_transfer_src_bit_arm = u64(0x00000004)
pub const tensor_usage_transfer_dst_bit_arm = u64(0x00000008)
pub const tensor_usage_image_aliasing_bit_arm = u64(0x00000010)
pub const tensor_usage_data_graph_bit_arm = u64(0x00000020)

// TensorDescriptionARM extends VkDataGraphPipelineResourceInfoARM,VkDataGraphPipelineConstantARM
pub type TensorDescriptionARM = C.VkTensorDescriptionARM

@[typedef]
pub struct C.VkTensorDescriptionARM {
pub mut:
	sType          StructureType = StructureType.tensor_description_arm
	pNext          voidptr       = unsafe { nil }
	tiling         TensorTilingARM
	format         Format
	dimensionCount u32
	pDimensions    &i64
	pStrides       &i64
	usage          TensorUsageFlagsARM
}

pub type TensorCreateInfoARM = C.VkTensorCreateInfoARM

@[typedef]
pub struct C.VkTensorCreateInfoARM {
pub mut:
	sType                 StructureType = StructureType.tensor_create_info_arm
	pNext                 voidptr       = unsafe { nil }
	flags                 TensorCreateFlagsARM
	pDescription          &TensorDescriptionARM
	sharingMode           SharingMode
	queueFamilyIndexCount u32
	pQueueFamilyIndices   &u32
}

pub type TensorViewCreateInfoARM = C.VkTensorViewCreateInfoARM

@[typedef]
pub struct C.VkTensorViewCreateInfoARM {
pub mut:
	sType  StructureType = StructureType.tensor_view_create_info_arm
	pNext  voidptr       = unsafe { nil }
	flags  TensorViewCreateFlagsARM
	tensor TensorARM
	format Format
}

pub type TensorMemoryRequirementsInfoARM = C.VkTensorMemoryRequirementsInfoARM

@[typedef]
pub struct C.VkTensorMemoryRequirementsInfoARM {
pub mut:
	sType  StructureType = StructureType.tensor_memory_requirements_info_arm
	pNext  voidptr       = unsafe { nil }
	tensor TensorARM
}

pub type BindTensorMemoryInfoARM = C.VkBindTensorMemoryInfoARM

@[typedef]
pub struct C.VkBindTensorMemoryInfoARM {
pub mut:
	sType        StructureType = StructureType.bind_tensor_memory_info_arm
	pNext        voidptr       = unsafe { nil }
	tensor       TensorARM
	memory       DeviceMemory
	memoryOffset DeviceSize
}

// WriteDescriptorSetTensorARM extends VkWriteDescriptorSet
pub type WriteDescriptorSetTensorARM = C.VkWriteDescriptorSetTensorARM

@[typedef]
pub struct C.VkWriteDescriptorSetTensorARM {
pub mut:
	sType           StructureType = StructureType.write_descriptor_set_tensor_arm
	pNext           voidptr       = unsafe { nil }
	tensorViewCount u32
	pTensorViews    &TensorViewARM
}

// TensorFormatPropertiesARM extends VkFormatProperties2
pub type TensorFormatPropertiesARM = C.VkTensorFormatPropertiesARM

@[typedef]
pub struct C.VkTensorFormatPropertiesARM {
pub mut:
	sType                       StructureType = StructureType.tensor_format_properties_arm
	pNext                       voidptr       = unsafe { nil }
	optimalTilingTensorFeatures FormatFeatureFlags2
	linearTilingTensorFeatures  FormatFeatureFlags2
}

// PhysicalDeviceTensorPropertiesARM extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceTensorPropertiesARM = C.VkPhysicalDeviceTensorPropertiesARM

@[typedef]
pub struct C.VkPhysicalDeviceTensorPropertiesARM {
pub mut:
	sType                                              StructureType = StructureType.physical_device_tensor_properties_arm
	pNext                                              voidptr       = unsafe { nil }
	maxTensorDimensionCount                            u32
	maxTensorElements                                  u64
	maxPerDimensionTensorElements                      u64
	maxTensorStride                                    i64
	maxTensorSize                                      u64
	maxTensorShaderAccessArrayLength                   u32
	maxTensorShaderAccessSize                          u32
	maxDescriptorSetStorageTensors                     u32
	maxPerStageDescriptorSetStorageTensors             u32
	maxDescriptorSetUpdateAfterBindStorageTensors      u32
	maxPerStageDescriptorUpdateAfterBindStorageTensors u32
	shaderStorageTensorArrayNonUniformIndexingNative   Bool32
	shaderTensorSupportedStages                        ShaderStageFlags
}

// TensorMemoryBarrierARM extends VkDependencyInfo
pub type TensorMemoryBarrierARM = C.VkTensorMemoryBarrierARM

@[typedef]
pub struct C.VkTensorMemoryBarrierARM {
pub mut:
	sType               StructureType = StructureType.tensor_memory_barrier_arm
	pNext               voidptr       = unsafe { nil }
	srcStageMask        PipelineStageFlags2
	srcAccessMask       AccessFlags2
	dstStageMask        PipelineStageFlags2
	dstAccessMask       AccessFlags2
	srcQueueFamilyIndex u32
	dstQueueFamilyIndex u32
	tensor              TensorARM
}

// TensorDependencyInfoARM extends VkDependencyInfo
pub type TensorDependencyInfoARM = C.VkTensorDependencyInfoARM

@[typedef]
pub struct C.VkTensorDependencyInfoARM {
pub mut:
	sType                    StructureType = StructureType.tensor_dependency_info_arm
	pNext                    voidptr       = unsafe { nil }
	tensorMemoryBarrierCount u32
	pTensorMemoryBarriers    &TensorMemoryBarrierARM
}

// PhysicalDeviceTensorFeaturesARM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceTensorFeaturesARM = C.VkPhysicalDeviceTensorFeaturesARM

@[typedef]
pub struct C.VkPhysicalDeviceTensorFeaturesARM {
pub mut:
	sType                                         StructureType = StructureType.physical_device_tensor_features_arm
	pNext                                         voidptr       = unsafe { nil }
	tensorNonPacked                               Bool32
	shaderTensorAccess                            Bool32
	shaderStorageTensorArrayDynamicIndexing       Bool32
	shaderStorageTensorArrayNonUniformIndexing    Bool32
	descriptorBindingStorageTensorUpdateAfterBind Bool32
	tensors                                       Bool32
}

pub type DeviceTensorMemoryRequirementsARM = C.VkDeviceTensorMemoryRequirementsARM

@[typedef]
pub struct C.VkDeviceTensorMemoryRequirementsARM {
pub mut:
	sType       StructureType = StructureType.device_tensor_memory_requirements_arm
	pNext       voidptr       = unsafe { nil }
	pCreateInfo &TensorCreateInfoARM
}

pub type TensorCopyARM = C.VkTensorCopyARM

@[typedef]
pub struct C.VkTensorCopyARM {
pub mut:
	sType          StructureType = StructureType.tensor_copy_arm
	pNext          voidptr       = unsafe { nil }
	dimensionCount u32
	pSrcOffset     &u64
	pDstOffset     &u64
	pExtent        &u64
}

pub type CopyTensorInfoARM = C.VkCopyTensorInfoARM

@[typedef]
pub struct C.VkCopyTensorInfoARM {
pub mut:
	sType       StructureType = StructureType.copy_tensor_info_arm
	pNext       voidptr       = unsafe { nil }
	srcTensor   TensorARM
	dstTensor   TensorARM
	regionCount u32
	pRegions    &TensorCopyARM
}

// MemoryDedicatedAllocateInfoTensorARM extends VkMemoryAllocateInfo
pub type MemoryDedicatedAllocateInfoTensorARM = C.VkMemoryDedicatedAllocateInfoTensorARM

@[typedef]
pub struct C.VkMemoryDedicatedAllocateInfoTensorARM {
pub mut:
	sType  StructureType = StructureType.memory_dedicated_allocate_info_tensor_arm
	pNext  voidptr       = unsafe { nil }
	tensor TensorARM
}

pub type PhysicalDeviceExternalTensorInfoARM = C.VkPhysicalDeviceExternalTensorInfoARM

@[typedef]
pub struct C.VkPhysicalDeviceExternalTensorInfoARM {
pub mut:
	sType        StructureType = StructureType.physical_device_external_tensor_info_arm
	pNext        voidptr       = unsafe { nil }
	flags        TensorCreateFlagsARM
	pDescription &TensorDescriptionARM
	handleType   ExternalMemoryHandleTypeFlagBits
}

pub type ExternalTensorPropertiesARM = C.VkExternalTensorPropertiesARM

@[typedef]
pub struct C.VkExternalTensorPropertiesARM {
pub mut:
	sType                    StructureType = StructureType.external_tensor_properties_arm
	pNext                    voidptr       = unsafe { nil }
	externalMemoryProperties ExternalMemoryProperties
}

// ExternalMemoryTensorCreateInfoARM extends VkTensorCreateInfoARM
pub type ExternalMemoryTensorCreateInfoARM = C.VkExternalMemoryTensorCreateInfoARM

@[typedef]
pub struct C.VkExternalMemoryTensorCreateInfoARM {
pub mut:
	sType       StructureType = StructureType.external_memory_tensor_create_info_arm
	pNext       voidptr       = unsafe { nil }
	handleTypes ExternalMemoryHandleTypeFlags
}

// PhysicalDeviceDescriptorBufferTensorFeaturesARM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDescriptorBufferTensorFeaturesARM = C.VkPhysicalDeviceDescriptorBufferTensorFeaturesARM

@[typedef]
pub struct C.VkPhysicalDeviceDescriptorBufferTensorFeaturesARM {
pub mut:
	sType                             StructureType = StructureType.physical_device_descriptor_buffer_tensor_features_arm
	pNext                             voidptr       = unsafe { nil }
	descriptorBufferTensorDescriptors Bool32
}

// PhysicalDeviceDescriptorBufferTensorPropertiesARM extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceDescriptorBufferTensorPropertiesARM = C.VkPhysicalDeviceDescriptorBufferTensorPropertiesARM

@[typedef]
pub struct C.VkPhysicalDeviceDescriptorBufferTensorPropertiesARM {
pub mut:
	sType                                     StructureType = StructureType.physical_device_descriptor_buffer_tensor_properties_arm
	pNext                                     voidptr       = unsafe { nil }
	tensorCaptureReplayDescriptorDataSize     usize
	tensorViewCaptureReplayDescriptorDataSize usize
	tensorDescriptorSize                      usize
}

// DescriptorGetTensorInfoARM extends VkDescriptorGetInfoEXT
pub type DescriptorGetTensorInfoARM = C.VkDescriptorGetTensorInfoARM

@[typedef]
pub struct C.VkDescriptorGetTensorInfoARM {
pub mut:
	sType      StructureType = StructureType.descriptor_get_tensor_info_arm
	pNext      voidptr       = unsafe { nil }
	tensorView TensorViewARM
}

pub type TensorCaptureDescriptorDataInfoARM = C.VkTensorCaptureDescriptorDataInfoARM

@[typedef]
pub struct C.VkTensorCaptureDescriptorDataInfoARM {
pub mut:
	sType  StructureType = StructureType.tensor_capture_descriptor_data_info_arm
	pNext  voidptr       = unsafe { nil }
	tensor TensorARM
}

pub type TensorViewCaptureDescriptorDataInfoARM = C.VkTensorViewCaptureDescriptorDataInfoARM

@[typedef]
pub struct C.VkTensorViewCaptureDescriptorDataInfoARM {
pub mut:
	sType      StructureType = StructureType.tensor_view_capture_descriptor_data_info_arm
	pNext      voidptr       = unsafe { nil }
	tensorView TensorViewARM
}

// FrameBoundaryTensorsARM extends VkSubmitInfo,VkSubmitInfo2,VkPresentInfoKHR,VkBindSparseInfo
pub type FrameBoundaryTensorsARM = C.VkFrameBoundaryTensorsARM

@[typedef]
pub struct C.VkFrameBoundaryTensorsARM {
pub mut:
	sType       StructureType = StructureType.frame_boundary_tensors_arm
	pNext       voidptr       = unsafe { nil }
	tensorCount u32
	pTensors    &TensorARM
}

@[keep_args_alive]
fn C.vkCreateTensorARM(device Device, p_create_info &TensorCreateInfoARM, p_allocator &AllocationCallbacks, p_tensor &TensorARM) Result

pub type PFN_vkCreateTensorARM = fn (device Device, p_create_info &TensorCreateInfoARM, p_allocator &AllocationCallbacks, p_tensor &TensorARM) Result

@[inline]
pub fn create_tensor_arm(device Device,
	p_create_info &TensorCreateInfoARM,
	p_allocator &AllocationCallbacks,
	p_tensor &TensorARM) Result {
	return C.vkCreateTensorARM(device, p_create_info, p_allocator, p_tensor)
}

@[keep_args_alive]
fn C.vkDestroyTensorARM(device Device, tensor TensorARM, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyTensorARM = fn (device Device, tensor TensorARM, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_tensor_arm(device Device,
	tensor TensorARM,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyTensorARM(device, tensor, p_allocator)
}

@[keep_args_alive]
fn C.vkCreateTensorViewARM(device Device, p_create_info &TensorViewCreateInfoARM, p_allocator &AllocationCallbacks, p_view &TensorViewARM) Result

pub type PFN_vkCreateTensorViewARM = fn (device Device, p_create_info &TensorViewCreateInfoARM, p_allocator &AllocationCallbacks, p_view &TensorViewARM) Result

@[inline]
pub fn create_tensor_view_arm(device Device,
	p_create_info &TensorViewCreateInfoARM,
	p_allocator &AllocationCallbacks,
	p_view &TensorViewARM) Result {
	return C.vkCreateTensorViewARM(device, p_create_info, p_allocator, p_view)
}

@[keep_args_alive]
fn C.vkDestroyTensorViewARM(device Device, tensor_view TensorViewARM, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyTensorViewARM = fn (device Device, tensor_view TensorViewARM, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_tensor_view_arm(device Device,
	tensor_view TensorViewARM,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyTensorViewARM(device, tensor_view, p_allocator)
}

@[keep_args_alive]
fn C.vkGetTensorMemoryRequirementsARM(device Device, p_info &TensorMemoryRequirementsInfoARM, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetTensorMemoryRequirementsARM = fn (device Device, p_info &TensorMemoryRequirementsInfoARM, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_tensor_memory_requirements_arm(device Device,
	p_info &TensorMemoryRequirementsInfoARM,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetTensorMemoryRequirementsARM(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkBindTensorMemoryARM(device Device, bind_info_count u32, p_bind_infos &BindTensorMemoryInfoARM) Result

pub type PFN_vkBindTensorMemoryARM = fn (device Device, bind_info_count u32, p_bind_infos &BindTensorMemoryInfoARM) Result

@[inline]
pub fn bind_tensor_memory_arm(device Device,
	bind_info_count u32,
	p_bind_infos &BindTensorMemoryInfoARM) Result {
	return C.vkBindTensorMemoryARM(device, bind_info_count, p_bind_infos)
}

@[keep_args_alive]
fn C.vkGetDeviceTensorMemoryRequirementsARM(device Device, p_info &DeviceTensorMemoryRequirementsARM, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetDeviceTensorMemoryRequirementsARM = fn (device Device, p_info &DeviceTensorMemoryRequirementsARM, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_device_tensor_memory_requirements_arm(device Device,
	p_info &DeviceTensorMemoryRequirementsARM,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetDeviceTensorMemoryRequirementsARM(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkCmdCopyTensorARM(command_buffer CommandBuffer, p_copy_tensor_info &CopyTensorInfoARM)

pub type PFN_vkCmdCopyTensorARM = fn (command_buffer CommandBuffer, p_copy_tensor_info &CopyTensorInfoARM)

@[inline]
pub fn cmd_copy_tensor_arm(command_buffer CommandBuffer,
	p_copy_tensor_info &CopyTensorInfoARM) {
	C.vkCmdCopyTensorARM(command_buffer, p_copy_tensor_info)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceExternalTensorPropertiesARM(physical_device PhysicalDevice, p_external_tensor_info &PhysicalDeviceExternalTensorInfoARM, mut p_external_tensor_properties ExternalTensorPropertiesARM)

pub type PFN_vkGetPhysicalDeviceExternalTensorPropertiesARM = fn (physical_device PhysicalDevice, p_external_tensor_info &PhysicalDeviceExternalTensorInfoARM, mut p_external_tensor_properties ExternalTensorPropertiesARM)

@[inline]
pub fn get_physical_device_external_tensor_properties_arm(physical_device PhysicalDevice,
	p_external_tensor_info &PhysicalDeviceExternalTensorInfoARM,
	mut p_external_tensor_properties ExternalTensorPropertiesARM) {
	C.vkGetPhysicalDeviceExternalTensorPropertiesARM(physical_device, p_external_tensor_info, mut
		p_external_tensor_properties)
}

@[keep_args_alive]
fn C.vkGetTensorOpaqueCaptureDescriptorDataARM(device Device, p_info &TensorCaptureDescriptorDataInfoARM, p_data voidptr) Result

pub type PFN_vkGetTensorOpaqueCaptureDescriptorDataARM = fn (device Device, p_info &TensorCaptureDescriptorDataInfoARM, p_data voidptr) Result

@[inline]
pub fn get_tensor_opaque_capture_descriptor_data_arm(device Device,
	p_info &TensorCaptureDescriptorDataInfoARM,
	p_data voidptr) Result {
	return C.vkGetTensorOpaqueCaptureDescriptorDataARM(device, p_info, p_data)
}

@[keep_args_alive]
fn C.vkGetTensorViewOpaqueCaptureDescriptorDataARM(device Device, p_info &TensorViewCaptureDescriptorDataInfoARM, p_data voidptr) Result

pub type PFN_vkGetTensorViewOpaqueCaptureDescriptorDataARM = fn (device Device, p_info &TensorViewCaptureDescriptorDataInfoARM, p_data voidptr) Result

@[inline]
pub fn get_tensor_view_opaque_capture_descriptor_data_arm(device Device,
	p_info &TensorViewCaptureDescriptorDataInfoARM,
	p_data voidptr) Result {
	return C.vkGetTensorViewOpaqueCaptureDescriptorDataARM(device, p_info, p_data)
}

pub const max_shader_module_identifier_size_ext = u32(32)
pub const ext_shader_module_identifier_spec_version = 1
pub const ext_shader_module_identifier_extension_name = c'VK_EXT_shader_module_identifier'
// PhysicalDeviceShaderModuleIdentifierFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderModuleIdentifierFeaturesEXT = C.VkPhysicalDeviceShaderModuleIdentifierFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderModuleIdentifierFeaturesEXT {
pub mut:
	sType                  StructureType = StructureType.physical_device_shader_module_identifier_features_ext
	pNext                  voidptr       = unsafe { nil }
	shaderModuleIdentifier Bool32
}

// PhysicalDeviceShaderModuleIdentifierPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceShaderModuleIdentifierPropertiesEXT = C.VkPhysicalDeviceShaderModuleIdentifierPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderModuleIdentifierPropertiesEXT {
pub mut:
	sType                               StructureType = StructureType.physical_device_shader_module_identifier_properties_ext
	pNext                               voidptr       = unsafe { nil }
	shaderModuleIdentifierAlgorithmUUID [uuid_size]u8
}

// PipelineShaderStageModuleIdentifierCreateInfoEXT extends VkPipelineShaderStageCreateInfo
pub type PipelineShaderStageModuleIdentifierCreateInfoEXT = C.VkPipelineShaderStageModuleIdentifierCreateInfoEXT

@[typedef]
pub struct C.VkPipelineShaderStageModuleIdentifierCreateInfoEXT {
pub mut:
	sType          StructureType = StructureType.pipeline_shader_stage_module_identifier_create_info_ext
	pNext          voidptr       = unsafe { nil }
	identifierSize u32
	pIdentifier    &u8
}

pub type ShaderModuleIdentifierEXT = C.VkShaderModuleIdentifierEXT

@[typedef]
pub struct C.VkShaderModuleIdentifierEXT {
pub mut:
	sType          StructureType = StructureType.shader_module_identifier_ext
	pNext          voidptr       = unsafe { nil }
	identifierSize u32
	identifier     [max_shader_module_identifier_size_ext]u8
}

@[keep_args_alive]
fn C.vkGetShaderModuleIdentifierEXT(device Device, shader_module ShaderModule, mut p_identifier ShaderModuleIdentifierEXT)

pub type PFN_vkGetShaderModuleIdentifierEXT = fn (device Device, shader_module ShaderModule, mut p_identifier ShaderModuleIdentifierEXT)

@[inline]
pub fn get_shader_module_identifier_ext(device Device,
	shader_module ShaderModule,
	mut p_identifier ShaderModuleIdentifierEXT) {
	C.vkGetShaderModuleIdentifierEXT(device, shader_module, mut p_identifier)
}

@[keep_args_alive]
fn C.vkGetShaderModuleCreateInfoIdentifierEXT(device Device, p_create_info &ShaderModuleCreateInfo, mut p_identifier ShaderModuleIdentifierEXT)

pub type PFN_vkGetShaderModuleCreateInfoIdentifierEXT = fn (device Device, p_create_info &ShaderModuleCreateInfo, mut p_identifier ShaderModuleIdentifierEXT)

@[inline]
pub fn get_shader_module_create_info_identifier_ext(device Device,
	p_create_info &ShaderModuleCreateInfo,
	mut p_identifier ShaderModuleIdentifierEXT) {
	C.vkGetShaderModuleCreateInfoIdentifierEXT(device, p_create_info, mut p_identifier)
}

pub const ext_rasterization_order_attachment_access_spec_version = 1
pub const ext_rasterization_order_attachment_access_extension_name = c'VK_EXT_rasterization_order_attachment_access'

// Pointer to VkOpticalFlowSessionNV_T
pub type OpticalFlowSessionNV = voidptr

pub const nv_optical_flow_spec_version = 1
pub const nv_optical_flow_extension_name = c'VK_NV_optical_flow'

pub enum OpticalFlowPerformanceLevelNV as u32 {
	unknown     = 0
	slow        = 1
	medium      = 2
	fast        = 3
	max_enum_nv = max_int
}

pub enum OpticalFlowSessionBindingPointNV as u32 {
	unknown              = 0
	input                = 1
	reference            = 2
	hint                 = 3
	flow_vector          = 4
	backward_flow_vector = 5
	cost                 = 6
	backward_cost        = 7
	global_flow          = 8
	max_enum_nv          = max_int
}

pub enum OpticalFlowGridSizeFlagBitsNV as u32 {
	unknown     = 0
	_1x1        = u32(0x00000001)
	_2x2        = u32(0x00000002)
	_4x4        = u32(0x00000004)
	_8x8        = u32(0x00000008)
	max_enum_nv = max_int
}
pub type OpticalFlowGridSizeFlagsNV = u32

pub enum OpticalFlowUsageFlagBitsNV as u32 {
	unknown     = 0
	input       = u32(0x00000001)
	output      = u32(0x00000002)
	hint        = u32(0x00000004)
	cost        = u32(0x00000008)
	global_flow = u32(0x00000010)
	max_enum_nv = max_int
}
pub type OpticalFlowUsageFlagsNV = u32

pub enum OpticalFlowSessionCreateFlagBitsNV as u32 {
	enable_hint        = u32(0x00000001)
	enable_cost        = u32(0x00000002)
	enable_global_flow = u32(0x00000004)
	allow_regions      = u32(0x00000008)
	both_directions    = u32(0x00000010)
	max_enum_nv        = max_int
}
pub type OpticalFlowSessionCreateFlagsNV = u32

pub enum OpticalFlowExecuteFlagBitsNV as u32 {
	disable_temporal_hints = u32(0x00000001)
	max_enum_nv            = max_int
}
pub type OpticalFlowExecuteFlagsNV = u32

// PhysicalDeviceOpticalFlowFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceOpticalFlowFeaturesNV = C.VkPhysicalDeviceOpticalFlowFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceOpticalFlowFeaturesNV {
pub mut:
	sType       StructureType = StructureType.physical_device_optical_flow_features_nv
	pNext       voidptr       = unsafe { nil }
	opticalFlow Bool32
}

// PhysicalDeviceOpticalFlowPropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceOpticalFlowPropertiesNV = C.VkPhysicalDeviceOpticalFlowPropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceOpticalFlowPropertiesNV {
pub mut:
	sType                      StructureType = StructureType.physical_device_optical_flow_properties_nv
	pNext                      voidptr       = unsafe { nil }
	supportedOutputGridSizes   OpticalFlowGridSizeFlagsNV
	supportedHintGridSizes     OpticalFlowGridSizeFlagsNV
	hintSupported              Bool32
	costSupported              Bool32
	bidirectionalFlowSupported Bool32
	globalFlowSupported        Bool32
	minWidth                   u32
	minHeight                  u32
	maxWidth                   u32
	maxHeight                  u32
	maxNumRegionsOfInterest    u32
}

// OpticalFlowImageFormatInfoNV extends VkPhysicalDeviceImageFormatInfo2,VkImageCreateInfo
pub type OpticalFlowImageFormatInfoNV = C.VkOpticalFlowImageFormatInfoNV

@[typedef]
pub struct C.VkOpticalFlowImageFormatInfoNV {
pub mut:
	sType StructureType = StructureType.optical_flow_image_format_info_nv
	pNext voidptr       = unsafe { nil }
	usage OpticalFlowUsageFlagsNV
}

pub type OpticalFlowImageFormatPropertiesNV = C.VkOpticalFlowImageFormatPropertiesNV

@[typedef]
pub struct C.VkOpticalFlowImageFormatPropertiesNV {
pub mut:
	sType  StructureType = StructureType.optical_flow_image_format_properties_nv
	pNext  voidptr       = unsafe { nil }
	format Format
}

pub type OpticalFlowSessionCreateInfoNV = C.VkOpticalFlowSessionCreateInfoNV

@[typedef]
pub struct C.VkOpticalFlowSessionCreateInfoNV {
pub mut:
	sType            StructureType = StructureType.optical_flow_session_create_info_nv
	pNext            voidptr       = unsafe { nil }
	width            u32
	height           u32
	imageFormat      Format
	flowVectorFormat Format
	costFormat       Format
	outputGridSize   OpticalFlowGridSizeFlagsNV
	hintGridSize     OpticalFlowGridSizeFlagsNV
	performanceLevel OpticalFlowPerformanceLevelNV
	flags            OpticalFlowSessionCreateFlagsNV
}

// OpticalFlowSessionCreatePrivateDataInfoNV extends VkOpticalFlowSessionCreateInfoNV
pub type OpticalFlowSessionCreatePrivateDataInfoNV = C.VkOpticalFlowSessionCreatePrivateDataInfoNV

@[typedef]
pub struct C.VkOpticalFlowSessionCreatePrivateDataInfoNV {
pub mut:
	sType        StructureType = StructureType.optical_flow_session_create_private_data_info_nv
	pNext        voidptr       = unsafe { nil }
	id           u32
	size         u32
	pPrivateData voidptr
}

pub type OpticalFlowExecuteInfoNV = C.VkOpticalFlowExecuteInfoNV

@[typedef]
pub struct C.VkOpticalFlowExecuteInfoNV {
pub mut:
	sType       StructureType = StructureType.optical_flow_execute_info_nv
	pNext       voidptr       = unsafe { nil }
	flags       OpticalFlowExecuteFlagsNV
	regionCount u32
	pRegions    &Rect2D
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceOpticalFlowImageFormatsNV(physical_device PhysicalDevice, p_optical_flow_image_format_info &OpticalFlowImageFormatInfoNV, p_format_count &u32, mut p_image_format_properties OpticalFlowImageFormatPropertiesNV) Result

pub type PFN_vkGetPhysicalDeviceOpticalFlowImageFormatsNV = fn (physical_device PhysicalDevice, p_optical_flow_image_format_info &OpticalFlowImageFormatInfoNV, p_format_count &u32, mut p_image_format_properties OpticalFlowImageFormatPropertiesNV) Result

@[inline]
pub fn get_physical_device_optical_flow_image_formats_nv(physical_device PhysicalDevice,
	p_optical_flow_image_format_info &OpticalFlowImageFormatInfoNV,
	p_format_count &u32,
	mut p_image_format_properties OpticalFlowImageFormatPropertiesNV) Result {
	return C.vkGetPhysicalDeviceOpticalFlowImageFormatsNV(physical_device, p_optical_flow_image_format_info,
		p_format_count, mut p_image_format_properties)
}

@[keep_args_alive]
fn C.vkCreateOpticalFlowSessionNV(device Device, p_create_info &OpticalFlowSessionCreateInfoNV, p_allocator &AllocationCallbacks, p_session &OpticalFlowSessionNV) Result

pub type PFN_vkCreateOpticalFlowSessionNV = fn (device Device, p_create_info &OpticalFlowSessionCreateInfoNV, p_allocator &AllocationCallbacks, p_session &OpticalFlowSessionNV) Result

@[inline]
pub fn create_optical_flow_session_nv(device Device,
	p_create_info &OpticalFlowSessionCreateInfoNV,
	p_allocator &AllocationCallbacks,
	p_session &OpticalFlowSessionNV) Result {
	return C.vkCreateOpticalFlowSessionNV(device, p_create_info, p_allocator, p_session)
}

@[keep_args_alive]
fn C.vkDestroyOpticalFlowSessionNV(device Device, session OpticalFlowSessionNV, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyOpticalFlowSessionNV = fn (device Device, session OpticalFlowSessionNV, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_optical_flow_session_nv(device Device,
	session OpticalFlowSessionNV,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyOpticalFlowSessionNV(device, session, p_allocator)
}

@[keep_args_alive]
fn C.vkBindOpticalFlowSessionImageNV(device Device, session OpticalFlowSessionNV, binding_point OpticalFlowSessionBindingPointNV, view ImageView, layout ImageLayout) Result

pub type PFN_vkBindOpticalFlowSessionImageNV = fn (device Device, session OpticalFlowSessionNV, binding_point OpticalFlowSessionBindingPointNV, view ImageView, layout ImageLayout) Result

@[inline]
pub fn bind_optical_flow_session_image_nv(device Device,
	session OpticalFlowSessionNV,
	binding_point OpticalFlowSessionBindingPointNV,
	view ImageView,
	layout ImageLayout) Result {
	return C.vkBindOpticalFlowSessionImageNV(device, session, binding_point, view, layout)
}

@[keep_args_alive]
fn C.vkCmdOpticalFlowExecuteNV(command_buffer CommandBuffer, session OpticalFlowSessionNV, p_execute_info &OpticalFlowExecuteInfoNV)

pub type PFN_vkCmdOpticalFlowExecuteNV = fn (command_buffer CommandBuffer, session OpticalFlowSessionNV, p_execute_info &OpticalFlowExecuteInfoNV)

@[inline]
pub fn cmd_optical_flow_execute_nv(command_buffer CommandBuffer,
	session OpticalFlowSessionNV,
	p_execute_info &OpticalFlowExecuteInfoNV) {
	C.vkCmdOpticalFlowExecuteNV(command_buffer, session, p_execute_info)
}

pub const ext_legacy_dithering_spec_version = 2
pub const ext_legacy_dithering_extension_name = c'VK_EXT_legacy_dithering'
// PhysicalDeviceLegacyDitheringFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceLegacyDitheringFeaturesEXT = C.VkPhysicalDeviceLegacyDitheringFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceLegacyDitheringFeaturesEXT {
pub mut:
	sType           StructureType = StructureType.physical_device_legacy_dithering_features_ext
	pNext           voidptr       = unsafe { nil }
	legacyDithering Bool32
}

pub const ext_pipeline_protected_access_spec_version = 1
pub const ext_pipeline_protected_access_extension_name = c'VK_EXT_pipeline_protected_access'

pub type PhysicalDevicePipelineProtectedAccessFeaturesEXT = C.VkPhysicalDevicePipelineProtectedAccessFeatures

pub const amd_anti_lag_spec_version = 1
pub const amd_anti_lag_extension_name = c'VK_AMD_anti_lag'

pub enum AntiLagModeAMD as u32 {
	driver_control = 0
	on             = 1
	off            = 2
	max_enum_amd   = max_int
}

pub enum AntiLagStageAMD as u32 {
	input        = 0
	present      = 1
	max_enum_amd = max_int
}
// PhysicalDeviceAntiLagFeaturesAMD extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceAntiLagFeaturesAMD = C.VkPhysicalDeviceAntiLagFeaturesAMD

@[typedef]
pub struct C.VkPhysicalDeviceAntiLagFeaturesAMD {
pub mut:
	sType   StructureType = StructureType.physical_device_anti_lag_features_amd
	pNext   voidptr       = unsafe { nil }
	antiLag Bool32
}

pub type AntiLagPresentationInfoAMD = C.VkAntiLagPresentationInfoAMD

@[typedef]
pub struct C.VkAntiLagPresentationInfoAMD {
pub mut:
	sType      StructureType = StructureType.anti_lag_presentation_info_amd
	pNext      voidptr       = unsafe { nil }
	stage      AntiLagStageAMD
	frameIndex u64
}

pub type AntiLagDataAMD = C.VkAntiLagDataAMD

@[typedef]
pub struct C.VkAntiLagDataAMD {
pub mut:
	sType             StructureType = StructureType.anti_lag_data_amd
	pNext             voidptr       = unsafe { nil }
	mode              AntiLagModeAMD
	maxFPS            u32
	pPresentationInfo &AntiLagPresentationInfoAMD
}

@[keep_args_alive]
fn C.vkAntiLagUpdateAMD(device Device, p_data &AntiLagDataAMD)

pub type PFN_vkAntiLagUpdateAMD = fn (device Device, p_data &AntiLagDataAMD)

@[inline]
pub fn anti_lag_update_amd(device Device,
	p_data &AntiLagDataAMD) {
	C.vkAntiLagUpdateAMD(device, p_data)
}

pub const amdx_dense_geometry_format_spec_version = 1
pub const amdx_dense_geometry_format_extension_name = c'VK_AMDX_dense_geometry_format'
pub const compressed_triangle_format_dgf1_byte_alignment_amdx = u32(128)
pub const compressed_triangle_format_dgf1_byte_stride_amdx = u32(128)

pub enum CompressedTriangleFormatAMDX as u32 {
	dgf1          = 0
	max_enum_amdx = max_int
}
// PhysicalDeviceDenseGeometryFormatFeaturesAMDX extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDenseGeometryFormatFeaturesAMDX = C.VkPhysicalDeviceDenseGeometryFormatFeaturesAMDX

@[typedef]
pub struct C.VkPhysicalDeviceDenseGeometryFormatFeaturesAMDX {
pub mut:
	sType               StructureType
	pNext               voidptr = unsafe { nil }
	denseGeometryFormat Bool32
}

// AccelerationStructureDenseGeometryFormatTrianglesDataAMDX extends VkAccelerationStructureGeometryKHR
pub type AccelerationStructureDenseGeometryFormatTrianglesDataAMDX = C.VkAccelerationStructureDenseGeometryFormatTrianglesDataAMDX

@[typedef]
pub struct C.VkAccelerationStructureDenseGeometryFormatTrianglesDataAMDX {
pub mut:
	sType             StructureType
	pNext             voidptr = unsafe { nil }
	compressedData    DeviceOrHostAddressConstKHR
	dataSize          DeviceSize
	numTriangles      u32
	numVertices       u32
	maxPrimitiveIndex u32
	maxGeometryIndex  u32
	format            CompressedTriangleFormatAMDX
}

// Pointer to VkShaderEXT_T
pub type ShaderEXT = voidptr

pub const ext_shader_object_spec_version = 1
pub const ext_shader_object_extension_name = c'VK_EXT_shader_object'

pub enum ShaderCodeTypeEXT as u32 {
	binary       = 0
	spirv        = 1
	max_enum_ext = max_int
}

pub enum DepthClampModeEXT as u32 {
	viewport_range     = 0
	user_defined_range = 1
	max_enum_ext       = max_int
}

pub enum ShaderCreateFlagBitsEXT as u32 {
	link_stage                       = u32(0x00000001)
	allow_varying_subgroup_size      = u32(0x00000002)
	require_full_subgroups           = u32(0x00000004)
	no_task_shader                   = u32(0x00000008)
	dispatch_base                    = u32(0x00000010)
	fragment_shading_rate_attachment = u32(0x00000020)
	fragment_density_map_attachment  = u32(0x00000040)
	indirect_bindable                = u32(0x00000080)
	_64_bit_indexing                 = u32(0x00008000)
	max_enum_ext                     = max_int
}
pub type ShaderCreateFlagsEXT = u32

// PhysicalDeviceShaderObjectFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderObjectFeaturesEXT = C.VkPhysicalDeviceShaderObjectFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderObjectFeaturesEXT {
pub mut:
	sType        StructureType = StructureType.physical_device_shader_object_features_ext
	pNext        voidptr       = unsafe { nil }
	shaderObject Bool32
}

// PhysicalDeviceShaderObjectPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceShaderObjectPropertiesEXT = C.VkPhysicalDeviceShaderObjectPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderObjectPropertiesEXT {
pub mut:
	sType               StructureType = StructureType.physical_device_shader_object_properties_ext
	pNext               voidptr       = unsafe { nil }
	shaderBinaryUUID    [uuid_size]u8
	shaderBinaryVersion u32
}

pub type ShaderCreateInfoEXT = C.VkShaderCreateInfoEXT

@[typedef]
pub struct C.VkShaderCreateInfoEXT {
pub mut:
	sType                  StructureType = StructureType.shader_create_info_ext
	pNext                  voidptr       = unsafe { nil }
	flags                  ShaderCreateFlagsEXT
	stage                  ShaderStageFlagBits
	nextStage              ShaderStageFlags
	codeType               ShaderCodeTypeEXT
	codeSize               usize
	pCode                  voidptr
	pName                  &char
	setLayoutCount         u32
	pSetLayouts            &DescriptorSetLayout
	pushConstantRangeCount u32
	pPushConstantRanges    &PushConstantRange
	pSpecializationInfo    &SpecializationInfo
}

pub type ShaderRequiredSubgroupSizeCreateInfoEXT = C.VkPipelineShaderStageRequiredSubgroupSizeCreateInfo

pub type DepthClampRangeEXT = C.VkDepthClampRangeEXT

@[typedef]
pub struct C.VkDepthClampRangeEXT {
pub mut:
	minDepthClamp f32
	maxDepthClamp f32
}

@[keep_args_alive]
fn C.vkCreateShadersEXT(device Device, create_info_count u32, p_create_infos &ShaderCreateInfoEXT, p_allocator &AllocationCallbacks, p_shaders &ShaderEXT) Result

pub type PFN_vkCreateShadersEXT = fn (device Device, create_info_count u32, p_create_infos &ShaderCreateInfoEXT, p_allocator &AllocationCallbacks, p_shaders &ShaderEXT) Result

@[inline]
pub fn create_shaders_ext(device Device,
	create_info_count u32,
	p_create_infos &ShaderCreateInfoEXT,
	p_allocator &AllocationCallbacks,
	p_shaders &ShaderEXT) Result {
	return C.vkCreateShadersEXT(device, create_info_count, p_create_infos, p_allocator,
		p_shaders)
}

@[keep_args_alive]
fn C.vkDestroyShaderEXT(device Device, shader ShaderEXT, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyShaderEXT = fn (device Device, shader ShaderEXT, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_shader_ext(device Device,
	shader ShaderEXT,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyShaderEXT(device, shader, p_allocator)
}

@[keep_args_alive]
fn C.vkGetShaderBinaryDataEXT(device Device, shader ShaderEXT, p_data_size &usize, p_data voidptr) Result

pub type PFN_vkGetShaderBinaryDataEXT = fn (device Device, shader ShaderEXT, p_data_size &usize, p_data voidptr) Result

@[inline]
pub fn get_shader_binary_data_ext(device Device,
	shader ShaderEXT,
	p_data_size &usize,
	p_data voidptr) Result {
	return C.vkGetShaderBinaryDataEXT(device, shader, p_data_size, p_data)
}

@[keep_args_alive]
fn C.vkCmdBindShadersEXT(command_buffer CommandBuffer, stage_count u32, p_stages &ShaderStageFlagBits, p_shaders &ShaderEXT)

pub type PFN_vkCmdBindShadersEXT = fn (command_buffer CommandBuffer, stage_count u32, p_stages &ShaderStageFlagBits, p_shaders &ShaderEXT)

@[inline]
pub fn cmd_bind_shaders_ext(command_buffer CommandBuffer,
	stage_count u32,
	p_stages &ShaderStageFlagBits,
	p_shaders &ShaderEXT) {
	C.vkCmdBindShadersEXT(command_buffer, stage_count, p_stages, p_shaders)
}

@[keep_args_alive]
fn C.vkCmdSetDepthClampRangeEXT(command_buffer CommandBuffer, depth_clamp_mode DepthClampModeEXT, p_depth_clamp_range &DepthClampRangeEXT)

pub type PFN_vkCmdSetDepthClampRangeEXT = fn (command_buffer CommandBuffer, depth_clamp_mode DepthClampModeEXT, p_depth_clamp_range &DepthClampRangeEXT)

@[inline]
pub fn cmd_set_depth_clamp_range_ext(command_buffer CommandBuffer,
	depth_clamp_mode DepthClampModeEXT,
	p_depth_clamp_range &DepthClampRangeEXT) {
	C.vkCmdSetDepthClampRangeEXT(command_buffer, depth_clamp_mode, p_depth_clamp_range)
}

pub const qcom_tile_properties_spec_version = 1
pub const qcom_tile_properties_extension_name = c'VK_QCOM_tile_properties'
// PhysicalDeviceTilePropertiesFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceTilePropertiesFeaturesQCOM = C.VkPhysicalDeviceTilePropertiesFeaturesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceTilePropertiesFeaturesQCOM {
pub mut:
	sType          StructureType = StructureType.physical_device_tile_properties_features_qcom
	pNext          voidptr       = unsafe { nil }
	tileProperties Bool32
}

pub type TilePropertiesQCOM = C.VkTilePropertiesQCOM

@[typedef]
pub struct C.VkTilePropertiesQCOM {
pub mut:
	sType     StructureType = StructureType.tile_properties_qcom
	pNext     voidptr       = unsafe { nil }
	tileSize  Extent3D
	apronSize Extent2D
	origin    Offset2D
}

@[keep_args_alive]
fn C.vkGetFramebufferTilePropertiesQCOM(device Device, framebuffer Framebuffer, p_properties_count &u32, mut p_properties TilePropertiesQCOM) Result

pub type PFN_vkGetFramebufferTilePropertiesQCOM = fn (device Device, framebuffer Framebuffer, p_properties_count &u32, mut p_properties TilePropertiesQCOM) Result

@[inline]
pub fn get_framebuffer_tile_properties_qcom(device Device,
	framebuffer Framebuffer,
	p_properties_count &u32,
	mut p_properties TilePropertiesQCOM) Result {
	return C.vkGetFramebufferTilePropertiesQCOM(device, framebuffer, p_properties_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkGetDynamicRenderingTilePropertiesQCOM(device Device, p_rendering_info &RenderingInfo, mut p_properties TilePropertiesQCOM) Result

pub type PFN_vkGetDynamicRenderingTilePropertiesQCOM = fn (device Device, p_rendering_info &RenderingInfo, mut p_properties TilePropertiesQCOM) Result

@[inline]
pub fn get_dynamic_rendering_tile_properties_qcom(device Device,
	p_rendering_info &RenderingInfo,
	mut p_properties TilePropertiesQCOM) Result {
	return C.vkGetDynamicRenderingTilePropertiesQCOM(device, p_rendering_info, mut p_properties)
}

pub const sec_amigo_profiling_spec_version = 1
pub const sec_amigo_profiling_extension_name = c'VK_SEC_amigo_profiling'
// PhysicalDeviceAmigoProfilingFeaturesSEC extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceAmigoProfilingFeaturesSEC = C.VkPhysicalDeviceAmigoProfilingFeaturesSEC

@[typedef]
pub struct C.VkPhysicalDeviceAmigoProfilingFeaturesSEC {
pub mut:
	sType          StructureType = StructureType.physical_device_amigo_profiling_features_sec
	pNext          voidptr       = unsafe { nil }
	amigoProfiling Bool32
}

// AmigoProfilingSubmitInfoSEC extends VkSubmitInfo
pub type AmigoProfilingSubmitInfoSEC = C.VkAmigoProfilingSubmitInfoSEC

@[typedef]
pub struct C.VkAmigoProfilingSubmitInfoSEC {
pub mut:
	sType               StructureType = StructureType.amigo_profiling_submit_info_sec
	pNext               voidptr       = unsafe { nil }
	firstDrawTimestamp  u64
	swapBufferTimestamp u64
}

pub const qcom_multiview_per_view_viewports_spec_version = 1
pub const qcom_multiview_per_view_viewports_extension_name = c'VK_QCOM_multiview_per_view_viewports'
// PhysicalDeviceMultiviewPerViewViewportsFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMultiviewPerViewViewportsFeaturesQCOM = C.VkPhysicalDeviceMultiviewPerViewViewportsFeaturesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceMultiviewPerViewViewportsFeaturesQCOM {
pub mut:
	sType                     StructureType = StructureType.physical_device_multiview_per_view_viewports_features_qcom
	pNext                     voidptr       = unsafe { nil }
	multiviewPerViewViewports Bool32
}

pub const nv_ray_tracing_invocation_reorder_spec_version = 1
pub const nv_ray_tracing_invocation_reorder_extension_name = c'VK_NV_ray_tracing_invocation_reorder'

pub enum RayTracingInvocationReorderModeNV as u32 {
	none        = 0
	reorder     = 1
	max_enum_nv = max_int
}
// PhysicalDeviceRayTracingInvocationReorderPropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceRayTracingInvocationReorderPropertiesNV = C.VkPhysicalDeviceRayTracingInvocationReorderPropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceRayTracingInvocationReorderPropertiesNV {
pub mut:
	sType                                     StructureType = StructureType.physical_device_ray_tracing_invocation_reorder_properties_nv
	pNext                                     voidptr       = unsafe { nil }
	rayTracingInvocationReorderReorderingHint RayTracingInvocationReorderModeNV
}

// PhysicalDeviceRayTracingInvocationReorderFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRayTracingInvocationReorderFeaturesNV = C.VkPhysicalDeviceRayTracingInvocationReorderFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceRayTracingInvocationReorderFeaturesNV {
pub mut:
	sType                       StructureType = StructureType.physical_device_ray_tracing_invocation_reorder_features_nv
	pNext                       voidptr       = unsafe { nil }
	rayTracingInvocationReorder Bool32
}

pub const nv_cooperative_vector_spec_version = 4
pub const nv_cooperative_vector_extension_name = c'VK_NV_cooperative_vector'

pub enum CooperativeVectorMatrixLayoutNV as u32 {
	row_major           = 0
	column_major        = 1
	inferencing_optimal = 2
	training_optimal    = 3
	max_enum_nv         = max_int
}
// PhysicalDeviceCooperativeVectorPropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceCooperativeVectorPropertiesNV = C.VkPhysicalDeviceCooperativeVectorPropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceCooperativeVectorPropertiesNV {
pub mut:
	sType                                        StructureType = StructureType.physical_device_cooperative_vector_properties_nv
	pNext                                        voidptr       = unsafe { nil }
	cooperativeVectorSupportedStages             ShaderStageFlags
	cooperativeVectorTrainingFloat16Accumulation Bool32
	cooperativeVectorTrainingFloat32Accumulation Bool32
	maxCooperativeVectorComponents               u32
}

// PhysicalDeviceCooperativeVectorFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCooperativeVectorFeaturesNV = C.VkPhysicalDeviceCooperativeVectorFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceCooperativeVectorFeaturesNV {
pub mut:
	sType                     StructureType = StructureType.physical_device_cooperative_vector_features_nv
	pNext                     voidptr       = unsafe { nil }
	cooperativeVector         Bool32
	cooperativeVectorTraining Bool32
}

pub type CooperativeVectorPropertiesNV = C.VkCooperativeVectorPropertiesNV

@[typedef]
pub struct C.VkCooperativeVectorPropertiesNV {
pub mut:
	sType                StructureType = StructureType.cooperative_vector_properties_nv
	pNext                voidptr       = unsafe { nil }
	inputType            ComponentTypeKHR
	inputInterpretation  ComponentTypeKHR
	matrixInterpretation ComponentTypeKHR
	biasInterpretation   ComponentTypeKHR
	resultType           ComponentTypeKHR
	transpose            Bool32
}

pub type ConvertCooperativeVectorMatrixInfoNV = C.VkConvertCooperativeVectorMatrixInfoNV

@[typedef]
pub struct C.VkConvertCooperativeVectorMatrixInfoNV {
pub mut:
	sType            StructureType = StructureType.convert_cooperative_vector_matrix_info_nv
	pNext            voidptr       = unsafe { nil }
	srcSize          usize
	srcData          DeviceOrHostAddressConstKHR
	pDstSize         &usize
	dstData          DeviceOrHostAddressKHR
	srcComponentType ComponentTypeKHR
	dstComponentType ComponentTypeKHR
	numRows          u32
	numColumns       u32
	srcLayout        CooperativeVectorMatrixLayoutNV
	srcStride        usize
	dstLayout        CooperativeVectorMatrixLayoutNV
	dstStride        usize
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceCooperativeVectorPropertiesNV(physical_device PhysicalDevice, p_property_count &u32, mut p_properties CooperativeVectorPropertiesNV) Result

pub type PFN_vkGetPhysicalDeviceCooperativeVectorPropertiesNV = fn (physical_device PhysicalDevice, p_property_count &u32, mut p_properties CooperativeVectorPropertiesNV) Result

@[inline]
pub fn get_physical_device_cooperative_vector_properties_nv(physical_device PhysicalDevice,
	p_property_count &u32,
	mut p_properties CooperativeVectorPropertiesNV) Result {
	return C.vkGetPhysicalDeviceCooperativeVectorPropertiesNV(physical_device, p_property_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkConvertCooperativeVectorMatrixNV(device Device, p_info &ConvertCooperativeVectorMatrixInfoNV) Result

pub type PFN_vkConvertCooperativeVectorMatrixNV = fn (device Device, p_info &ConvertCooperativeVectorMatrixInfoNV) Result

@[inline]
pub fn convert_cooperative_vector_matrix_nv(device Device,
	p_info &ConvertCooperativeVectorMatrixInfoNV) Result {
	return C.vkConvertCooperativeVectorMatrixNV(device, p_info)
}

@[keep_args_alive]
fn C.vkCmdConvertCooperativeVectorMatrixNV(command_buffer CommandBuffer, info_count u32, p_infos &ConvertCooperativeVectorMatrixInfoNV)

pub type PFN_vkCmdConvertCooperativeVectorMatrixNV = fn (command_buffer CommandBuffer, info_count u32, p_infos &ConvertCooperativeVectorMatrixInfoNV)

@[inline]
pub fn cmd_convert_cooperative_vector_matrix_nv(command_buffer CommandBuffer,
	info_count u32,
	p_infos &ConvertCooperativeVectorMatrixInfoNV) {
	C.vkCmdConvertCooperativeVectorMatrixNV(command_buffer, info_count, p_infos)
}

pub const nv_extended_sparse_address_space_spec_version = 1
pub const nv_extended_sparse_address_space_extension_name = c'VK_NV_extended_sparse_address_space'
// PhysicalDeviceExtendedSparseAddressSpaceFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceExtendedSparseAddressSpaceFeaturesNV = C.VkPhysicalDeviceExtendedSparseAddressSpaceFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceExtendedSparseAddressSpaceFeaturesNV {
pub mut:
	sType                      StructureType = StructureType.physical_device_extended_sparse_address_space_features_nv
	pNext                      voidptr       = unsafe { nil }
	extendedSparseAddressSpace Bool32
}

// PhysicalDeviceExtendedSparseAddressSpacePropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceExtendedSparseAddressSpacePropertiesNV = C.VkPhysicalDeviceExtendedSparseAddressSpacePropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceExtendedSparseAddressSpacePropertiesNV {
pub mut:
	sType                          StructureType = StructureType.physical_device_extended_sparse_address_space_properties_nv
	pNext                          voidptr       = unsafe { nil }
	extendedSparseAddressSpaceSize DeviceSize
	extendedSparseImageUsageFlags  ImageUsageFlags
	extendedSparseBufferUsageFlags BufferUsageFlags
}

pub const ext_mutable_descriptor_type_spec_version = 1
pub const ext_mutable_descriptor_type_extension_name = c'VK_EXT_mutable_descriptor_type'

pub const ext_legacy_vertex_attributes_spec_version = 1
pub const ext_legacy_vertex_attributes_extension_name = c'VK_EXT_legacy_vertex_attributes'
// PhysicalDeviceLegacyVertexAttributesFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceLegacyVertexAttributesFeaturesEXT = C.VkPhysicalDeviceLegacyVertexAttributesFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceLegacyVertexAttributesFeaturesEXT {
pub mut:
	sType                  StructureType = StructureType.physical_device_legacy_vertex_attributes_features_ext
	pNext                  voidptr       = unsafe { nil }
	legacyVertexAttributes Bool32
}

// PhysicalDeviceLegacyVertexAttributesPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceLegacyVertexAttributesPropertiesEXT = C.VkPhysicalDeviceLegacyVertexAttributesPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceLegacyVertexAttributesPropertiesEXT {
pub mut:
	sType                      StructureType = StructureType.physical_device_legacy_vertex_attributes_properties_ext
	pNext                      voidptr       = unsafe { nil }
	nativeUnalignedPerformance Bool32
}

pub const ext_layer_settings_spec_version = 2
pub const ext_layer_settings_extension_name = c'VK_EXT_layer_settings'

pub enum LayerSettingTypeEXT as u32 {
	bool32       = 0
	int32        = 1
	int64        = 2
	uint32       = 3
	uint64       = 4
	float32      = 5
	float64      = 6
	string       = 7
	max_enum_ext = max_int
}
pub type LayerSettingEXT = C.VkLayerSettingEXT

@[typedef]
pub struct C.VkLayerSettingEXT {
pub mut:
	pLayerName   &char
	pSettingName &char
	type         LayerSettingTypeEXT
	valueCount   u32
	pValues      voidptr
}

// LayerSettingsCreateInfoEXT extends VkInstanceCreateInfo
pub type LayerSettingsCreateInfoEXT = C.VkLayerSettingsCreateInfoEXT

@[typedef]
pub struct C.VkLayerSettingsCreateInfoEXT {
pub mut:
	sType        StructureType = StructureType.layer_settings_create_info_ext
	pNext        voidptr       = unsafe { nil }
	settingCount u32
	pSettings    &LayerSettingEXT
}

pub const arm_shader_core_builtins_spec_version = 2
pub const arm_shader_core_builtins_extension_name = c'VK_ARM_shader_core_builtins'
// PhysicalDeviceShaderCoreBuiltinsFeaturesARM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderCoreBuiltinsFeaturesARM = C.VkPhysicalDeviceShaderCoreBuiltinsFeaturesARM

@[typedef]
pub struct C.VkPhysicalDeviceShaderCoreBuiltinsFeaturesARM {
pub mut:
	sType              StructureType = StructureType.physical_device_shader_core_builtins_features_arm
	pNext              voidptr       = unsafe { nil }
	shaderCoreBuiltins Bool32
}

// PhysicalDeviceShaderCoreBuiltinsPropertiesARM extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceShaderCoreBuiltinsPropertiesARM = C.VkPhysicalDeviceShaderCoreBuiltinsPropertiesARM

@[typedef]
pub struct C.VkPhysicalDeviceShaderCoreBuiltinsPropertiesARM {
pub mut:
	sType              StructureType = StructureType.physical_device_shader_core_builtins_properties_arm
	pNext              voidptr       = unsafe { nil }
	shaderCoreMask     u64
	shaderCoreCount    u32
	shaderWarpsPerCore u32
}

pub const ext_pipeline_library_group_handles_spec_version = 1
pub const ext_pipeline_library_group_handles_extension_name = c'VK_EXT_pipeline_library_group_handles'
// PhysicalDevicePipelineLibraryGroupHandlesFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePipelineLibraryGroupHandlesFeaturesEXT = C.VkPhysicalDevicePipelineLibraryGroupHandlesFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDevicePipelineLibraryGroupHandlesFeaturesEXT {
pub mut:
	sType                       StructureType = StructureType.physical_device_pipeline_library_group_handles_features_ext
	pNext                       voidptr       = unsafe { nil }
	pipelineLibraryGroupHandles Bool32
}

pub const ext_dynamic_rendering_unused_attachments_spec_version = 1
pub const ext_dynamic_rendering_unused_attachments_extension_name = c'VK_EXT_dynamic_rendering_unused_attachments'
// PhysicalDeviceDynamicRenderingUnusedAttachmentsFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDynamicRenderingUnusedAttachmentsFeaturesEXT = C.VkPhysicalDeviceDynamicRenderingUnusedAttachmentsFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDynamicRenderingUnusedAttachmentsFeaturesEXT {
pub mut:
	sType                             StructureType = StructureType.physical_device_dynamic_rendering_unused_attachments_features_ext
	pNext                             voidptr       = unsafe { nil }
	dynamicRenderingUnusedAttachments Bool32
}

pub const nv_low_latency_2_spec_version = 2
pub const nv_low_latency_2_extension_name = c'VK_NV_low_latency2'

pub enum LatencyMarkerNV as u32 {
	simulation_start               = 0
	simulation_end                 = 1
	rendersubmit_start             = 2
	rendersubmit_end               = 3
	present_start                  = 4
	present_end                    = 5
	input_sample                   = 6
	trigger_flash                  = 7
	out_of_band_rendersubmit_start = 8
	out_of_band_rendersubmit_end   = 9
	out_of_band_present_start      = 10
	out_of_band_present_end        = 11
	max_enum_nv                    = max_int
}

pub enum OutOfBandQueueTypeNV as u32 {
	render      = 0
	present     = 1
	max_enum_nv = max_int
}
pub type LatencySleepModeInfoNV = C.VkLatencySleepModeInfoNV

@[typedef]
pub struct C.VkLatencySleepModeInfoNV {
pub mut:
	sType             StructureType = StructureType.latency_sleep_mode_info_nv
	pNext             voidptr       = unsafe { nil }
	lowLatencyMode    Bool32
	lowLatencyBoost   Bool32
	minimumIntervalUs u32
}

pub type LatencySleepInfoNV = C.VkLatencySleepInfoNV

@[typedef]
pub struct C.VkLatencySleepInfoNV {
pub mut:
	sType           StructureType = StructureType.latency_sleep_info_nv
	pNext           voidptr       = unsafe { nil }
	signalSemaphore Semaphore
	value           u64
}

pub type SetLatencyMarkerInfoNV = C.VkSetLatencyMarkerInfoNV

@[typedef]
pub struct C.VkSetLatencyMarkerInfoNV {
pub mut:
	sType     StructureType = StructureType.set_latency_marker_info_nv
	pNext     voidptr       = unsafe { nil }
	presentID u64
	marker    LatencyMarkerNV
}

pub type LatencyTimingsFrameReportNV = C.VkLatencyTimingsFrameReportNV

@[typedef]
pub struct C.VkLatencyTimingsFrameReportNV {
pub mut:
	sType                    StructureType = StructureType.latency_timings_frame_report_nv
	pNext                    voidptr       = unsafe { nil }
	presentID                u64
	inputSampleTimeUs        u64
	simStartTimeUs           u64
	simEndTimeUs             u64
	renderSubmitStartTimeUs  u64
	renderSubmitEndTimeUs    u64
	presentStartTimeUs       u64
	presentEndTimeUs         u64
	driverStartTimeUs        u64
	driverEndTimeUs          u64
	osRenderQueueStartTimeUs u64
	osRenderQueueEndTimeUs   u64
	gpuRenderStartTimeUs     u64
	gpuRenderEndTimeUs       u64
}

pub type GetLatencyMarkerInfoNV = C.VkGetLatencyMarkerInfoNV

@[typedef]
pub struct C.VkGetLatencyMarkerInfoNV {
pub mut:
	sType       StructureType = StructureType.get_latency_marker_info_nv
	pNext       voidptr       = unsafe { nil }
	timingCount u32
	pTimings    &LatencyTimingsFrameReportNV
}

// LatencySubmissionPresentIdNV extends VkSubmitInfo,VkSubmitInfo2
pub type LatencySubmissionPresentIdNV = C.VkLatencySubmissionPresentIdNV

@[typedef]
pub struct C.VkLatencySubmissionPresentIdNV {
pub mut:
	sType     StructureType = StructureType.latency_submission_present_id_nv
	pNext     voidptr       = unsafe { nil }
	presentID u64
}

// SwapchainLatencyCreateInfoNV extends VkSwapchainCreateInfoKHR
pub type SwapchainLatencyCreateInfoNV = C.VkSwapchainLatencyCreateInfoNV

@[typedef]
pub struct C.VkSwapchainLatencyCreateInfoNV {
pub mut:
	sType             StructureType = StructureType.swapchain_latency_create_info_nv
	pNext             voidptr       = unsafe { nil }
	latencyModeEnable Bool32
}

pub type OutOfBandQueueTypeInfoNV = C.VkOutOfBandQueueTypeInfoNV

@[typedef]
pub struct C.VkOutOfBandQueueTypeInfoNV {
pub mut:
	sType     StructureType = StructureType.out_of_band_queue_type_info_nv
	pNext     voidptr       = unsafe { nil }
	queueType OutOfBandQueueTypeNV
}

// LatencySurfaceCapabilitiesNV extends VkSurfaceCapabilities2KHR
pub type LatencySurfaceCapabilitiesNV = C.VkLatencySurfaceCapabilitiesNV

@[typedef]
pub struct C.VkLatencySurfaceCapabilitiesNV {
pub mut:
	sType            StructureType = StructureType.latency_surface_capabilities_nv
	pNext            voidptr       = unsafe { nil }
	presentModeCount u32
	pPresentModes    &PresentModeKHR
}

@[keep_args_alive]
fn C.vkSetLatencySleepModeNV(device Device, swapchain SwapchainKHR, p_sleep_mode_info &LatencySleepModeInfoNV) Result

pub type PFN_vkSetLatencySleepModeNV = fn (device Device, swapchain SwapchainKHR, p_sleep_mode_info &LatencySleepModeInfoNV) Result

@[inline]
pub fn set_latency_sleep_mode_nv(device Device,
	swapchain SwapchainKHR,
	p_sleep_mode_info &LatencySleepModeInfoNV) Result {
	return C.vkSetLatencySleepModeNV(device, swapchain, p_sleep_mode_info)
}

@[keep_args_alive]
fn C.vkLatencySleepNV(device Device, swapchain SwapchainKHR, p_sleep_info &LatencySleepInfoNV) Result

pub type PFN_vkLatencySleepNV = fn (device Device, swapchain SwapchainKHR, p_sleep_info &LatencySleepInfoNV) Result

@[inline]
pub fn latency_sleep_nv(device Device,
	swapchain SwapchainKHR,
	p_sleep_info &LatencySleepInfoNV) Result {
	return C.vkLatencySleepNV(device, swapchain, p_sleep_info)
}

@[keep_args_alive]
fn C.vkSetLatencyMarkerNV(device Device, swapchain SwapchainKHR, p_latency_marker_info &SetLatencyMarkerInfoNV)

pub type PFN_vkSetLatencyMarkerNV = fn (device Device, swapchain SwapchainKHR, p_latency_marker_info &SetLatencyMarkerInfoNV)

@[inline]
pub fn set_latency_marker_nv(device Device,
	swapchain SwapchainKHR,
	p_latency_marker_info &SetLatencyMarkerInfoNV) {
	C.vkSetLatencyMarkerNV(device, swapchain, p_latency_marker_info)
}

@[keep_args_alive]
fn C.vkGetLatencyTimingsNV(device Device, swapchain SwapchainKHR, mut p_latency_marker_info GetLatencyMarkerInfoNV)

pub type PFN_vkGetLatencyTimingsNV = fn (device Device, swapchain SwapchainKHR, mut p_latency_marker_info GetLatencyMarkerInfoNV)

@[inline]
pub fn get_latency_timings_nv(device Device,
	swapchain SwapchainKHR,
	mut p_latency_marker_info GetLatencyMarkerInfoNV) {
	C.vkGetLatencyTimingsNV(device, swapchain, mut p_latency_marker_info)
}

@[keep_args_alive]
fn C.vkQueueNotifyOutOfBandNV(queue Queue, p_queue_type_info &OutOfBandQueueTypeInfoNV)

pub type PFN_vkQueueNotifyOutOfBandNV = fn (queue Queue, p_queue_type_info &OutOfBandQueueTypeInfoNV)

@[inline]
pub fn queue_notify_out_of_band_nv(queue Queue,
	p_queue_type_info &OutOfBandQueueTypeInfoNV) {
	C.vkQueueNotifyOutOfBandNV(queue, p_queue_type_info)
}

// Pointer to VkDataGraphPipelineSessionARM_T
pub type DataGraphPipelineSessionARM = voidptr

pub const max_physical_device_data_graph_operation_set_name_size_arm = u32(128)
pub const arm_data_graph_spec_version = 1
pub const arm_data_graph_extension_name = c'VK_ARM_data_graph'

pub enum DataGraphPipelineSessionBindPointARM as u32 {
	transient    = 0
	max_enum_arm = max_int
}

pub enum DataGraphPipelineSessionBindPointTypeARM as u32 {
	memory       = 0
	max_enum_arm = max_int
}

pub enum DataGraphPipelinePropertyARM as u32 {
	creation_log = 0
	identifier   = 1
	max_enum_arm = max_int
}

pub enum PhysicalDeviceDataGraphProcessingEngineTypeARM as u32 {
	default      = 0
	max_enum_arm = max_int
}

pub enum PhysicalDeviceDataGraphOperationTypeARM as u32 {
	spirv_extended_instruction_set = 0
	max_enum_arm                   = max_int
}
pub type DataGraphPipelineSessionCreateFlagsARM = u64

// Flag bits for DataGraphPipelineSessionCreateFlagBitsARM
pub type DataGraphPipelineSessionCreateFlagBitsARM = u64

pub const data_graph_pipeline_session_create_protected_bit_arm = u64(0x00000001)

pub type DataGraphPipelineDispatchFlagsARM = u64

// Flag bits for DataGraphPipelineDispatchFlagBitsARM
pub type DataGraphPipelineDispatchFlagBitsARM = u64

// PhysicalDeviceDataGraphFeaturesARM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDataGraphFeaturesARM = C.VkPhysicalDeviceDataGraphFeaturesARM

@[typedef]
pub struct C.VkPhysicalDeviceDataGraphFeaturesARM {
pub mut:
	sType                            StructureType = StructureType.physical_device_data_graph_features_arm
	pNext                            voidptr       = unsafe { nil }
	dataGraph                        Bool32
	dataGraphUpdateAfterBind         Bool32
	dataGraphSpecializationConstants Bool32
	dataGraphDescriptorBuffer        Bool32
	dataGraphShaderModule            Bool32
}

pub type DataGraphPipelineConstantARM = C.VkDataGraphPipelineConstantARM

@[typedef]
pub struct C.VkDataGraphPipelineConstantARM {
pub mut:
	sType         StructureType = StructureType.data_graph_pipeline_constant_arm
	pNext         voidptr       = unsafe { nil }
	id            u32
	pConstantData voidptr
}

pub type DataGraphPipelineResourceInfoARM = C.VkDataGraphPipelineResourceInfoARM

@[typedef]
pub struct C.VkDataGraphPipelineResourceInfoARM {
pub mut:
	sType         StructureType = StructureType.data_graph_pipeline_resource_info_arm
	pNext         voidptr       = unsafe { nil }
	descriptorSet u32
	binding       u32
	arrayElement  u32
}

// DataGraphPipelineCompilerControlCreateInfoARM extends VkDataGraphPipelineCreateInfoARM
pub type DataGraphPipelineCompilerControlCreateInfoARM = C.VkDataGraphPipelineCompilerControlCreateInfoARM

@[typedef]
pub struct C.VkDataGraphPipelineCompilerControlCreateInfoARM {
pub mut:
	sType          StructureType = StructureType.data_graph_pipeline_compiler_control_create_info_arm
	pNext          voidptr       = unsafe { nil }
	pVendorOptions &char
}

pub type DataGraphPipelineCreateInfoARM = C.VkDataGraphPipelineCreateInfoARM

@[typedef]
pub struct C.VkDataGraphPipelineCreateInfoARM {
pub mut:
	sType             StructureType = StructureType.data_graph_pipeline_create_info_arm
	pNext             voidptr       = unsafe { nil }
	flags             PipelineCreateFlags2KHR
	layout            PipelineLayout
	resourceInfoCount u32
	pResourceInfos    &DataGraphPipelineResourceInfoARM
}

// DataGraphPipelineShaderModuleCreateInfoARM extends VkDataGraphPipelineCreateInfoARM
pub type DataGraphPipelineShaderModuleCreateInfoARM = C.VkDataGraphPipelineShaderModuleCreateInfoARM

@[typedef]
pub struct C.VkDataGraphPipelineShaderModuleCreateInfoARM {
pub mut:
	sType               StructureType = StructureType.data_graph_pipeline_shader_module_create_info_arm
	pNext               voidptr       = unsafe { nil }
	module              ShaderModule
	pName               &char
	pSpecializationInfo &SpecializationInfo
	constantCount       u32
	pConstants          &DataGraphPipelineConstantARM
}

pub type DataGraphPipelineSessionCreateInfoARM = C.VkDataGraphPipelineSessionCreateInfoARM

@[typedef]
pub struct C.VkDataGraphPipelineSessionCreateInfoARM {
pub mut:
	sType             StructureType = StructureType.data_graph_pipeline_session_create_info_arm
	pNext             voidptr       = unsafe { nil }
	flags             DataGraphPipelineSessionCreateFlagsARM
	dataGraphPipeline Pipeline
}

pub type DataGraphPipelineSessionBindPointRequirementsInfoARM = C.VkDataGraphPipelineSessionBindPointRequirementsInfoARM

@[typedef]
pub struct C.VkDataGraphPipelineSessionBindPointRequirementsInfoARM {
pub mut:
	sType   StructureType = StructureType.data_graph_pipeline_session_bind_point_requirements_info_arm
	pNext   voidptr       = unsafe { nil }
	session DataGraphPipelineSessionARM
}

pub type DataGraphPipelineSessionBindPointRequirementARM = C.VkDataGraphPipelineSessionBindPointRequirementARM

@[typedef]
pub struct C.VkDataGraphPipelineSessionBindPointRequirementARM {
pub mut:
	sType         StructureType = StructureType.data_graph_pipeline_session_bind_point_requirement_arm
	pNext         voidptr       = unsafe { nil }
	bindPoint     DataGraphPipelineSessionBindPointARM
	bindPointType DataGraphPipelineSessionBindPointTypeARM
	numObjects    u32
}

pub type DataGraphPipelineSessionMemoryRequirementsInfoARM = C.VkDataGraphPipelineSessionMemoryRequirementsInfoARM

@[typedef]
pub struct C.VkDataGraphPipelineSessionMemoryRequirementsInfoARM {
pub mut:
	sType       StructureType = StructureType.data_graph_pipeline_session_memory_requirements_info_arm
	pNext       voidptr       = unsafe { nil }
	session     DataGraphPipelineSessionARM
	bindPoint   DataGraphPipelineSessionBindPointARM
	objectIndex u32
}

pub type BindDataGraphPipelineSessionMemoryInfoARM = C.VkBindDataGraphPipelineSessionMemoryInfoARM

@[typedef]
pub struct C.VkBindDataGraphPipelineSessionMemoryInfoARM {
pub mut:
	sType        StructureType = StructureType.bind_data_graph_pipeline_session_memory_info_arm
	pNext        voidptr       = unsafe { nil }
	session      DataGraphPipelineSessionARM
	bindPoint    DataGraphPipelineSessionBindPointARM
	objectIndex  u32
	memory       DeviceMemory
	memoryOffset DeviceSize
}

pub type DataGraphPipelineInfoARM = C.VkDataGraphPipelineInfoARM

@[typedef]
pub struct C.VkDataGraphPipelineInfoARM {
pub mut:
	sType             StructureType = StructureType.data_graph_pipeline_info_arm
	pNext             voidptr       = unsafe { nil }
	dataGraphPipeline Pipeline
}

pub type DataGraphPipelinePropertyQueryResultARM = C.VkDataGraphPipelinePropertyQueryResultARM

@[typedef]
pub struct C.VkDataGraphPipelinePropertyQueryResultARM {
pub mut:
	sType    StructureType = StructureType.data_graph_pipeline_property_query_result_arm
	pNext    voidptr       = unsafe { nil }
	property DataGraphPipelinePropertyARM
	isText   Bool32
	dataSize usize
	pData    voidptr
}

// DataGraphPipelineIdentifierCreateInfoARM extends VkDataGraphPipelineCreateInfoARM
pub type DataGraphPipelineIdentifierCreateInfoARM = C.VkDataGraphPipelineIdentifierCreateInfoARM

@[typedef]
pub struct C.VkDataGraphPipelineIdentifierCreateInfoARM {
pub mut:
	sType          StructureType = StructureType.data_graph_pipeline_identifier_create_info_arm
	pNext          voidptr       = unsafe { nil }
	identifierSize u32
	pIdentifier    &u8
}

pub type DataGraphPipelineDispatchInfoARM = C.VkDataGraphPipelineDispatchInfoARM

@[typedef]
pub struct C.VkDataGraphPipelineDispatchInfoARM {
pub mut:
	sType StructureType = StructureType.data_graph_pipeline_dispatch_info_arm
	pNext voidptr       = unsafe { nil }
	flags DataGraphPipelineDispatchFlagsARM
}

pub type PhysicalDeviceDataGraphProcessingEngineARM = C.VkPhysicalDeviceDataGraphProcessingEngineARM

@[typedef]
pub struct C.VkPhysicalDeviceDataGraphProcessingEngineARM {
pub mut:
	type      PhysicalDeviceDataGraphProcessingEngineTypeARM
	isForeign Bool32
}

pub type PhysicalDeviceDataGraphOperationSupportARM = C.VkPhysicalDeviceDataGraphOperationSupportARM

@[typedef]
pub struct C.VkPhysicalDeviceDataGraphOperationSupportARM {
pub mut:
	operationType PhysicalDeviceDataGraphOperationTypeARM
	name          [max_physical_device_data_graph_operation_set_name_size_arm]char
	version       u32
}

pub type QueueFamilyDataGraphPropertiesARM = C.VkQueueFamilyDataGraphPropertiesARM

@[typedef]
pub struct C.VkQueueFamilyDataGraphPropertiesARM {
pub mut:
	sType     StructureType = StructureType.queue_family_data_graph_properties_arm
	pNext     voidptr       = unsafe { nil }
	engine    PhysicalDeviceDataGraphProcessingEngineARM
	operation PhysicalDeviceDataGraphOperationSupportARM
}

// DataGraphProcessingEngineCreateInfoARM extends VkDataGraphPipelineCreateInfoARM,VkDescriptorPoolCreateInfo,VkCommandPoolCreateInfo
pub type DataGraphProcessingEngineCreateInfoARM = C.VkDataGraphProcessingEngineCreateInfoARM

@[typedef]
pub struct C.VkDataGraphProcessingEngineCreateInfoARM {
pub mut:
	sType                 StructureType = StructureType.data_graph_processing_engine_create_info_arm
	pNext                 voidptr       = unsafe { nil }
	processingEngineCount u32
	pProcessingEngines    &PhysicalDeviceDataGraphProcessingEngineARM
}

pub type PhysicalDeviceQueueFamilyDataGraphProcessingEngineInfoARM = C.VkPhysicalDeviceQueueFamilyDataGraphProcessingEngineInfoARM

@[typedef]
pub struct C.VkPhysicalDeviceQueueFamilyDataGraphProcessingEngineInfoARM {
pub mut:
	sType            StructureType = StructureType.physical_device_queue_family_data_graph_processing_engine_info_arm
	pNext            voidptr       = unsafe { nil }
	queueFamilyIndex u32
	engineType       PhysicalDeviceDataGraphProcessingEngineTypeARM
}

pub type QueueFamilyDataGraphProcessingEnginePropertiesARM = C.VkQueueFamilyDataGraphProcessingEnginePropertiesARM

@[typedef]
pub struct C.VkQueueFamilyDataGraphProcessingEnginePropertiesARM {
pub mut:
	sType                       StructureType = StructureType.queue_family_data_graph_processing_engine_properties_arm
	pNext                       voidptr       = unsafe { nil }
	foreignSemaphoreHandleTypes ExternalSemaphoreHandleTypeFlags
	foreignMemoryHandleTypes    ExternalMemoryHandleTypeFlags
}

// DataGraphPipelineConstantTensorSemiStructuredSparsityInfoARM extends VkDataGraphPipelineConstantARM
pub type DataGraphPipelineConstantTensorSemiStructuredSparsityInfoARM = C.VkDataGraphPipelineConstantTensorSemiStructuredSparsityInfoARM

@[typedef]
pub struct C.VkDataGraphPipelineConstantTensorSemiStructuredSparsityInfoARM {
pub mut:
	sType     StructureType = StructureType.data_graph_pipeline_constant_tensor_semi_structured_sparsity_info_arm
	pNext     voidptr       = unsafe { nil }
	dimension u32
	zeroCount u32
	groupSize u32
}

@[keep_args_alive]
fn C.vkCreateDataGraphPipelinesARM(device Device, deferred_operation DeferredOperationKHR, pipeline_cache PipelineCache, create_info_count u32, p_create_infos &DataGraphPipelineCreateInfoARM, p_allocator &AllocationCallbacks, p_pipelines &Pipeline) Result

pub type PFN_vkCreateDataGraphPipelinesARM = fn (device Device, deferred_operation DeferredOperationKHR, pipeline_cache PipelineCache, create_info_count u32, p_create_infos &DataGraphPipelineCreateInfoARM, p_allocator &AllocationCallbacks, p_pipelines &Pipeline) Result

@[inline]
pub fn create_data_graph_pipelines_arm(device Device,
	deferred_operation DeferredOperationKHR,
	pipeline_cache PipelineCache,
	create_info_count u32,
	p_create_infos &DataGraphPipelineCreateInfoARM,
	p_allocator &AllocationCallbacks,
	p_pipelines &Pipeline) Result {
	return C.vkCreateDataGraphPipelinesARM(device, deferred_operation, pipeline_cache,
		create_info_count, p_create_infos, p_allocator, p_pipelines)
}

@[keep_args_alive]
fn C.vkCreateDataGraphPipelineSessionARM(device Device, p_create_info &DataGraphPipelineSessionCreateInfoARM, p_allocator &AllocationCallbacks, p_session &DataGraphPipelineSessionARM) Result

pub type PFN_vkCreateDataGraphPipelineSessionARM = fn (device Device, p_create_info &DataGraphPipelineSessionCreateInfoARM, p_allocator &AllocationCallbacks, p_session &DataGraphPipelineSessionARM) Result

@[inline]
pub fn create_data_graph_pipeline_session_arm(device Device,
	p_create_info &DataGraphPipelineSessionCreateInfoARM,
	p_allocator &AllocationCallbacks,
	p_session &DataGraphPipelineSessionARM) Result {
	return C.vkCreateDataGraphPipelineSessionARM(device, p_create_info, p_allocator, p_session)
}

@[keep_args_alive]
fn C.vkGetDataGraphPipelineSessionBindPointRequirementsARM(device Device, p_info &DataGraphPipelineSessionBindPointRequirementsInfoARM, p_bind_point_requirement_count &u32, mut p_bind_point_requirements DataGraphPipelineSessionBindPointRequirementARM) Result

pub type PFN_vkGetDataGraphPipelineSessionBindPointRequirementsARM = fn (device Device, p_info &DataGraphPipelineSessionBindPointRequirementsInfoARM, p_bind_point_requirement_count &u32, mut p_bind_point_requirements DataGraphPipelineSessionBindPointRequirementARM) Result

@[inline]
pub fn get_data_graph_pipeline_session_bind_point_requirements_arm(device Device,
	p_info &DataGraphPipelineSessionBindPointRequirementsInfoARM,
	p_bind_point_requirement_count &u32,
	mut p_bind_point_requirements DataGraphPipelineSessionBindPointRequirementARM) Result {
	return C.vkGetDataGraphPipelineSessionBindPointRequirementsARM(device, p_info, p_bind_point_requirement_count, mut
		p_bind_point_requirements)
}

@[keep_args_alive]
fn C.vkGetDataGraphPipelineSessionMemoryRequirementsARM(device Device, p_info &DataGraphPipelineSessionMemoryRequirementsInfoARM, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetDataGraphPipelineSessionMemoryRequirementsARM = fn (device Device, p_info &DataGraphPipelineSessionMemoryRequirementsInfoARM, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_data_graph_pipeline_session_memory_requirements_arm(device Device,
	p_info &DataGraphPipelineSessionMemoryRequirementsInfoARM,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetDataGraphPipelineSessionMemoryRequirementsARM(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkBindDataGraphPipelineSessionMemoryARM(device Device, bind_info_count u32, p_bind_infos &BindDataGraphPipelineSessionMemoryInfoARM) Result

pub type PFN_vkBindDataGraphPipelineSessionMemoryARM = fn (device Device, bind_info_count u32, p_bind_infos &BindDataGraphPipelineSessionMemoryInfoARM) Result

@[inline]
pub fn bind_data_graph_pipeline_session_memory_arm(device Device,
	bind_info_count u32,
	p_bind_infos &BindDataGraphPipelineSessionMemoryInfoARM) Result {
	return C.vkBindDataGraphPipelineSessionMemoryARM(device, bind_info_count, p_bind_infos)
}

@[keep_args_alive]
fn C.vkDestroyDataGraphPipelineSessionARM(device Device, session DataGraphPipelineSessionARM, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyDataGraphPipelineSessionARM = fn (device Device, session DataGraphPipelineSessionARM, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_data_graph_pipeline_session_arm(device Device,
	session DataGraphPipelineSessionARM,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyDataGraphPipelineSessionARM(device, session, p_allocator)
}

@[keep_args_alive]
fn C.vkCmdDispatchDataGraphARM(command_buffer CommandBuffer, session DataGraphPipelineSessionARM, p_info &DataGraphPipelineDispatchInfoARM)

pub type PFN_vkCmdDispatchDataGraphARM = fn (command_buffer CommandBuffer, session DataGraphPipelineSessionARM, p_info &DataGraphPipelineDispatchInfoARM)

@[inline]
pub fn cmd_dispatch_data_graph_arm(command_buffer CommandBuffer,
	session DataGraphPipelineSessionARM,
	p_info &DataGraphPipelineDispatchInfoARM) {
	C.vkCmdDispatchDataGraphARM(command_buffer, session, p_info)
}

@[keep_args_alive]
fn C.vkGetDataGraphPipelineAvailablePropertiesARM(device Device, p_pipeline_info &DataGraphPipelineInfoARM, p_properties_count &u32, p_properties &DataGraphPipelinePropertyARM) Result

pub type PFN_vkGetDataGraphPipelineAvailablePropertiesARM = fn (device Device, p_pipeline_info &DataGraphPipelineInfoARM, p_properties_count &u32, p_properties &DataGraphPipelinePropertyARM) Result

@[inline]
pub fn get_data_graph_pipeline_available_properties_arm(device Device,
	p_pipeline_info &DataGraphPipelineInfoARM,
	p_properties_count &u32,
	p_properties &DataGraphPipelinePropertyARM) Result {
	return C.vkGetDataGraphPipelineAvailablePropertiesARM(device, p_pipeline_info, p_properties_count,
		p_properties)
}

@[keep_args_alive]
fn C.vkGetDataGraphPipelinePropertiesARM(device Device, p_pipeline_info &DataGraphPipelineInfoARM, properties_count u32, mut p_properties DataGraphPipelinePropertyQueryResultARM) Result

pub type PFN_vkGetDataGraphPipelinePropertiesARM = fn (device Device, p_pipeline_info &DataGraphPipelineInfoARM, properties_count u32, mut p_properties DataGraphPipelinePropertyQueryResultARM) Result

@[inline]
pub fn get_data_graph_pipeline_properties_arm(device Device,
	p_pipeline_info &DataGraphPipelineInfoARM,
	properties_count u32,
	mut p_properties DataGraphPipelinePropertyQueryResultARM) Result {
	return C.vkGetDataGraphPipelinePropertiesARM(device, p_pipeline_info, properties_count, mut
		p_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceQueueFamilyDataGraphPropertiesARM(physical_device PhysicalDevice, queue_family_index u32, p_queue_family_data_graph_property_count &u32, mut p_queue_family_data_graph_properties QueueFamilyDataGraphPropertiesARM) Result

pub type PFN_vkGetPhysicalDeviceQueueFamilyDataGraphPropertiesARM = fn (physical_device PhysicalDevice, queue_family_index u32, p_queue_family_data_graph_property_count &u32, mut p_queue_family_data_graph_properties QueueFamilyDataGraphPropertiesARM) Result

@[inline]
pub fn get_physical_device_queue_family_data_graph_properties_arm(physical_device PhysicalDevice,
	queue_family_index u32,
	p_queue_family_data_graph_property_count &u32,
	mut p_queue_family_data_graph_properties QueueFamilyDataGraphPropertiesARM) Result {
	return C.vkGetPhysicalDeviceQueueFamilyDataGraphPropertiesARM(physical_device, queue_family_index,
		p_queue_family_data_graph_property_count, mut p_queue_family_data_graph_properties)
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceQueueFamilyDataGraphProcessingEnginePropertiesARM(physical_device PhysicalDevice, p_queue_family_data_graph_processing_engine_info &PhysicalDeviceQueueFamilyDataGraphProcessingEngineInfoARM, mut p_queue_family_data_graph_processing_engine_properties QueueFamilyDataGraphProcessingEnginePropertiesARM)

pub type PFN_vkGetPhysicalDeviceQueueFamilyDataGraphProcessingEnginePropertiesARM = fn (physical_device PhysicalDevice, p_queue_family_data_graph_processing_engine_info &PhysicalDeviceQueueFamilyDataGraphProcessingEngineInfoARM, mut p_queue_family_data_graph_processing_engine_properties QueueFamilyDataGraphProcessingEnginePropertiesARM)

@[inline]
pub fn get_physical_device_queue_family_data_graph_processing_engine_properties_arm(physical_device PhysicalDevice,
	p_queue_family_data_graph_processing_engine_info &PhysicalDeviceQueueFamilyDataGraphProcessingEngineInfoARM,
	mut p_queue_family_data_graph_processing_engine_properties QueueFamilyDataGraphProcessingEnginePropertiesARM) {
	C.vkGetPhysicalDeviceQueueFamilyDataGraphProcessingEnginePropertiesARM(physical_device,
		p_queue_family_data_graph_processing_engine_info, mut p_queue_family_data_graph_processing_engine_properties)
}

pub const qcom_multiview_per_view_render_areas_spec_version = 1
pub const qcom_multiview_per_view_render_areas_extension_name = c'VK_QCOM_multiview_per_view_render_areas'
// PhysicalDeviceMultiviewPerViewRenderAreasFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMultiviewPerViewRenderAreasFeaturesQCOM = C.VkPhysicalDeviceMultiviewPerViewRenderAreasFeaturesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceMultiviewPerViewRenderAreasFeaturesQCOM {
pub mut:
	sType                       StructureType = StructureType.physical_device_multiview_per_view_render_areas_features_qcom
	pNext                       voidptr       = unsafe { nil }
	multiviewPerViewRenderAreas Bool32
}

// MultiviewPerViewRenderAreasRenderPassBeginInfoQCOM extends VkRenderPassBeginInfo,VkRenderingInfo
pub type MultiviewPerViewRenderAreasRenderPassBeginInfoQCOM = C.VkMultiviewPerViewRenderAreasRenderPassBeginInfoQCOM

@[typedef]
pub struct C.VkMultiviewPerViewRenderAreasRenderPassBeginInfoQCOM {
pub mut:
	sType                  StructureType = StructureType.multiview_per_view_render_areas_render_pass_begin_info_qcom
	pNext                  voidptr       = unsafe { nil }
	perViewRenderAreaCount u32
	pPerViewRenderAreas    &Rect2D
}

pub const nv_per_stage_descriptor_set_spec_version = 1
pub const nv_per_stage_descriptor_set_extension_name = c'VK_NV_per_stage_descriptor_set'
// PhysicalDevicePerStageDescriptorSetFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePerStageDescriptorSetFeaturesNV = C.VkPhysicalDevicePerStageDescriptorSetFeaturesNV

@[typedef]
pub struct C.VkPhysicalDevicePerStageDescriptorSetFeaturesNV {
pub mut:
	sType                 StructureType = StructureType.physical_device_per_stage_descriptor_set_features_nv
	pNext                 voidptr       = unsafe { nil }
	perStageDescriptorSet Bool32
	dynamicPipelineLayout Bool32
}

pub const qcom_image_processing_2_spec_version = 1
pub const qcom_image_processing_2_extension_name = c'VK_QCOM_image_processing2'

pub enum BlockMatchWindowCompareModeQCOM as u32 {
	min           = 0
	max           = 1
	max_enum_qcom = max_int
}
// PhysicalDeviceImageProcessing2FeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceImageProcessing2FeaturesQCOM = C.VkPhysicalDeviceImageProcessing2FeaturesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceImageProcessing2FeaturesQCOM {
pub mut:
	sType              StructureType = StructureType.physical_device_image_processing2_features_qcom
	pNext              voidptr       = unsafe { nil }
	textureBlockMatch2 Bool32
}

// PhysicalDeviceImageProcessing2PropertiesQCOM extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceImageProcessing2PropertiesQCOM = C.VkPhysicalDeviceImageProcessing2PropertiesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceImageProcessing2PropertiesQCOM {
pub mut:
	sType               StructureType = StructureType.physical_device_image_processing2_properties_qcom
	pNext               voidptr       = unsafe { nil }
	maxBlockMatchWindow Extent2D
}

// SamplerBlockMatchWindowCreateInfoQCOM extends VkSamplerCreateInfo
pub type SamplerBlockMatchWindowCreateInfoQCOM = C.VkSamplerBlockMatchWindowCreateInfoQCOM

@[typedef]
pub struct C.VkSamplerBlockMatchWindowCreateInfoQCOM {
pub mut:
	sType             StructureType = StructureType.sampler_block_match_window_create_info_qcom
	pNext             voidptr       = unsafe { nil }
	windowExtent      Extent2D
	windowCompareMode BlockMatchWindowCompareModeQCOM
}

pub const qcom_filter_cubic_weights_spec_version = 1
pub const qcom_filter_cubic_weights_extension_name = c'VK_QCOM_filter_cubic_weights'

pub enum CubicFilterWeightsQCOM as u32 {
	catmull_rom           = 0
	zero_tangent_cardinal = 1
	b_spline              = 2
	mitchell_netravali    = 3
	max_enum_qcom         = max_int
}
// PhysicalDeviceCubicWeightsFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCubicWeightsFeaturesQCOM = C.VkPhysicalDeviceCubicWeightsFeaturesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceCubicWeightsFeaturesQCOM {
pub mut:
	sType                  StructureType = StructureType.physical_device_cubic_weights_features_qcom
	pNext                  voidptr       = unsafe { nil }
	selectableCubicWeights Bool32
}

// SamplerCubicWeightsCreateInfoQCOM extends VkSamplerCreateInfo
pub type SamplerCubicWeightsCreateInfoQCOM = C.VkSamplerCubicWeightsCreateInfoQCOM

@[typedef]
pub struct C.VkSamplerCubicWeightsCreateInfoQCOM {
pub mut:
	sType        StructureType = StructureType.sampler_cubic_weights_create_info_qcom
	pNext        voidptr       = unsafe { nil }
	cubicWeights CubicFilterWeightsQCOM
}

// BlitImageCubicWeightsInfoQCOM extends VkBlitImageInfo2
pub type BlitImageCubicWeightsInfoQCOM = C.VkBlitImageCubicWeightsInfoQCOM

@[typedef]
pub struct C.VkBlitImageCubicWeightsInfoQCOM {
pub mut:
	sType        StructureType = StructureType.blit_image_cubic_weights_info_qcom
	pNext        voidptr       = unsafe { nil }
	cubicWeights CubicFilterWeightsQCOM
}

pub const qcom_ycbcr_degamma_spec_version = 1
pub const qcom_ycbcr_degamma_extension_name = c'VK_QCOM_ycbcr_degamma'
// PhysicalDeviceYcbcrDegammaFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceYcbcrDegammaFeaturesQCOM = C.VkPhysicalDeviceYcbcrDegammaFeaturesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceYcbcrDegammaFeaturesQCOM {
pub mut:
	sType        StructureType = StructureType.physical_device_ycbcr_degamma_features_qcom
	pNext        voidptr       = unsafe { nil }
	ycbcrDegamma Bool32
}

// SamplerYcbcrConversionYcbcrDegammaCreateInfoQCOM extends VkSamplerYcbcrConversionCreateInfo
pub type SamplerYcbcrConversionYcbcrDegammaCreateInfoQCOM = C.VkSamplerYcbcrConversionYcbcrDegammaCreateInfoQCOM

@[typedef]
pub struct C.VkSamplerYcbcrConversionYcbcrDegammaCreateInfoQCOM {
pub mut:
	sType             StructureType = StructureType.sampler_ycbcr_conversion_ycbcr_degamma_create_info_qcom
	pNext             voidptr       = unsafe { nil }
	enableYDegamma    Bool32
	enableCbCrDegamma Bool32
}

pub const qcom_filter_cubic_clamp_spec_version = 1
pub const qcom_filter_cubic_clamp_extension_name = c'VK_QCOM_filter_cubic_clamp'
// PhysicalDeviceCubicClampFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCubicClampFeaturesQCOM = C.VkPhysicalDeviceCubicClampFeaturesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceCubicClampFeaturesQCOM {
pub mut:
	sType           StructureType = StructureType.physical_device_cubic_clamp_features_qcom
	pNext           voidptr       = unsafe { nil }
	cubicRangeClamp Bool32
}

pub const ext_attachment_feedback_loop_dynamic_state_spec_version = 1
pub const ext_attachment_feedback_loop_dynamic_state_extension_name = c'VK_EXT_attachment_feedback_loop_dynamic_state'
// PhysicalDeviceAttachmentFeedbackLoopDynamicStateFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceAttachmentFeedbackLoopDynamicStateFeaturesEXT = C.VkPhysicalDeviceAttachmentFeedbackLoopDynamicStateFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceAttachmentFeedbackLoopDynamicStateFeaturesEXT {
pub mut:
	sType                              StructureType = StructureType.physical_device_attachment_feedback_loop_dynamic_state_features_ext
	pNext                              voidptr       = unsafe { nil }
	attachmentFeedbackLoopDynamicState Bool32
}

@[keep_args_alive]
fn C.vkCmdSetAttachmentFeedbackLoopEnableEXT(command_buffer CommandBuffer, aspect_mask ImageAspectFlags)

pub type PFN_vkCmdSetAttachmentFeedbackLoopEnableEXT = fn (command_buffer CommandBuffer, aspect_mask ImageAspectFlags)

@[inline]
pub fn cmd_set_attachment_feedback_loop_enable_ext(command_buffer CommandBuffer,
	aspect_mask ImageAspectFlags) {
	C.vkCmdSetAttachmentFeedbackLoopEnableEXT(command_buffer, aspect_mask)
}

pub const msft_layered_driver_spec_version = 1
pub const msft_layered_driver_extension_name = c'VK_MST_layered_driver'

pub enum LayeredDriverUnderlyingApiMSFT as u32 {
	none          = 0
	d3d12         = 1
	max_enum_msft = max_int
}
// PhysicalDeviceLayeredDriverPropertiesMSFT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceLayeredDriverPropertiesMSFT = C.VkPhysicalDeviceLayeredDriverPropertiesMSFT

@[typedef]
pub struct C.VkPhysicalDeviceLayeredDriverPropertiesMSFT {
pub mut:
	sType         StructureType = StructureType.physical_device_layered_driver_properties_msft
	pNext         voidptr       = unsafe { nil }
	underlyingAPI LayeredDriverUnderlyingApiMSFT
}

pub const nv_descriptor_pool_overallocation_spec_version = 1
pub const nv_descriptor_pool_overallocation_extension_name = c'VK_NV_descriptor_pool_overallocation'
// PhysicalDeviceDescriptorPoolOverallocationFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDescriptorPoolOverallocationFeaturesNV = C.VkPhysicalDeviceDescriptorPoolOverallocationFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceDescriptorPoolOverallocationFeaturesNV {
pub mut:
	sType                        StructureType = StructureType.physical_device_descriptor_pool_overallocation_features_nv
	pNext                        voidptr       = unsafe { nil }
	descriptorPoolOverallocation Bool32
}

pub const qcom_tile_memory_heap_spec_version = 1
pub const qcom_tile_memory_heap_extension_name = c'VK_QCOM_tile_memory_heap'
// PhysicalDeviceTileMemoryHeapFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceTileMemoryHeapFeaturesQCOM = C.VkPhysicalDeviceTileMemoryHeapFeaturesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceTileMemoryHeapFeaturesQCOM {
pub mut:
	sType          StructureType = StructureType.physical_device_tile_memory_heap_features_qcom
	pNext          voidptr       = unsafe { nil }
	tileMemoryHeap Bool32
}

// PhysicalDeviceTileMemoryHeapPropertiesQCOM extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceTileMemoryHeapPropertiesQCOM = C.VkPhysicalDeviceTileMemoryHeapPropertiesQCOM

@[typedef]
pub struct C.VkPhysicalDeviceTileMemoryHeapPropertiesQCOM {
pub mut:
	sType               StructureType = StructureType.physical_device_tile_memory_heap_properties_qcom
	pNext               voidptr       = unsafe { nil }
	queueSubmitBoundary Bool32
	tileBufferTransfers Bool32
}

// TileMemoryRequirementsQCOM extends VkMemoryRequirements2
pub type TileMemoryRequirementsQCOM = C.VkTileMemoryRequirementsQCOM

@[typedef]
pub struct C.VkTileMemoryRequirementsQCOM {
pub mut:
	sType     StructureType = StructureType.tile_memory_requirements_qcom
	pNext     voidptr       = unsafe { nil }
	size      DeviceSize
	alignment DeviceSize
}

// TileMemoryBindInfoQCOM extends VkCommandBufferInheritanceInfo
pub type TileMemoryBindInfoQCOM = C.VkTileMemoryBindInfoQCOM

@[typedef]
pub struct C.VkTileMemoryBindInfoQCOM {
pub mut:
	sType  StructureType = StructureType.tile_memory_bind_info_qcom
	pNext  voidptr       = unsafe { nil }
	memory DeviceMemory
}

// TileMemorySizeInfoQCOM extends VkRenderPassCreateInfo,VkRenderPassCreateInfo2,VkRenderingInfo
pub type TileMemorySizeInfoQCOM = C.VkTileMemorySizeInfoQCOM

@[typedef]
pub struct C.VkTileMemorySizeInfoQCOM {
pub mut:
	sType StructureType = StructureType.tile_memory_size_info_qcom
	pNext voidptr       = unsafe { nil }
	size  DeviceSize
}

@[keep_args_alive]
fn C.vkCmdBindTileMemoryQCOM(command_buffer CommandBuffer, p_tile_memory_bind_info &TileMemoryBindInfoQCOM)

pub type PFN_vkCmdBindTileMemoryQCOM = fn (command_buffer CommandBuffer, p_tile_memory_bind_info &TileMemoryBindInfoQCOM)

@[inline]
pub fn cmd_bind_tile_memory_qcom(command_buffer CommandBuffer,
	p_tile_memory_bind_info &TileMemoryBindInfoQCOM) {
	C.vkCmdBindTileMemoryQCOM(command_buffer, p_tile_memory_bind_info)
}

pub const ext_memory_decompression_spec_version = 1
pub const ext_memory_decompression_extension_name = c'VK_EXT_memory_decompression'

pub type DecompressMemoryRegionEXT = C.VkDecompressMemoryRegionEXT

@[typedef]
pub struct C.VkDecompressMemoryRegionEXT {
pub mut:
	srcAddress       DeviceAddress
	dstAddress       DeviceAddress
	compressedSize   DeviceSize
	decompressedSize DeviceSize
}

pub type DecompressMemoryInfoEXT = C.VkDecompressMemoryInfoEXT

@[typedef]
pub struct C.VkDecompressMemoryInfoEXT {
pub mut:
	sType               StructureType = StructureType.decompress_memory_info_ext
	pNext               voidptr       = unsafe { nil }
	decompressionMethod MemoryDecompressionMethodFlagsEXT
	regionCount         u32
	pRegions            &DecompressMemoryRegionEXT
}

@[keep_args_alive]
fn C.vkCmdDecompressMemoryEXT(command_buffer CommandBuffer, p_decompress_memory_info_ext &DecompressMemoryInfoEXT)

pub type PFN_vkCmdDecompressMemoryEXT = fn (command_buffer CommandBuffer, p_decompress_memory_info_ext &DecompressMemoryInfoEXT)

@[inline]
pub fn cmd_decompress_memory_ext(command_buffer CommandBuffer,
	p_decompress_memory_info_ext &DecompressMemoryInfoEXT) {
	C.vkCmdDecompressMemoryEXT(command_buffer, p_decompress_memory_info_ext)
}

@[keep_args_alive]
fn C.vkCmdDecompressMemoryIndirectCountEXT(command_buffer CommandBuffer, decompression_method MemoryDecompressionMethodFlagsEXT, indirect_commands_address DeviceAddress, indirect_commands_count_address DeviceAddress, max_decompression_count u32, stride u32)

pub type PFN_vkCmdDecompressMemoryIndirectCountEXT = fn (command_buffer CommandBuffer, decompression_method MemoryDecompressionMethodFlagsEXT, indirect_commands_address DeviceAddress, indirect_commands_count_address DeviceAddress, max_decompression_count u32, stride u32)

@[inline]
pub fn cmd_decompress_memory_indirect_count_ext(command_buffer CommandBuffer,
	decompression_method MemoryDecompressionMethodFlagsEXT,
	indirect_commands_address DeviceAddress,
	indirect_commands_count_address DeviceAddress,
	max_decompression_count u32,
	stride u32) {
	C.vkCmdDecompressMemoryIndirectCountEXT(command_buffer, decompression_method, indirect_commands_address,
		indirect_commands_count_address, max_decompression_count, stride)
}

pub const nv_display_stereo_spec_version = 1
pub const nv_display_stereo_extension_name = c'VK_NV_display_stereo'

pub enum DisplaySurfaceStereoTypeNV as u32 {
	none               = 0
	onboard_din        = 1
	hdmi3d             = 2
	inband_displayport = 3
	max_enum_nv        = max_int
}
// DisplaySurfaceStereoCreateInfoNV extends VkDisplaySurfaceCreateInfoKHR
pub type DisplaySurfaceStereoCreateInfoNV = C.VkDisplaySurfaceStereoCreateInfoNV

@[typedef]
pub struct C.VkDisplaySurfaceStereoCreateInfoNV {
pub mut:
	sType      StructureType = StructureType.display_surface_stereo_create_info_nv
	pNext      voidptr       = unsafe { nil }
	stereoType DisplaySurfaceStereoTypeNV
}

// DisplayModeStereoPropertiesNV extends VkDisplayModeProperties2KHR
pub type DisplayModeStereoPropertiesNV = C.VkDisplayModeStereoPropertiesNV

@[typedef]
pub struct C.VkDisplayModeStereoPropertiesNV {
pub mut:
	sType           StructureType = StructureType.display_mode_stereo_properties_nv
	pNext           voidptr       = unsafe { nil }
	hdmi3DSupported Bool32
}

pub const nv_raw_access_chains_spec_version = 1
pub const nv_raw_access_chains_extension_name = c'VK_NV_raw_access_chains'
// PhysicalDeviceRawAccessChainsFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRawAccessChainsFeaturesNV = C.VkPhysicalDeviceRawAccessChainsFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceRawAccessChainsFeaturesNV {
pub mut:
	sType                 StructureType = StructureType.physical_device_raw_access_chains_features_nv
	pNext                 voidptr       = unsafe { nil }
	shaderRawAccessChains Bool32
}

// Pointer to VkExternalComputeQueueNV_T
pub type ExternalComputeQueueNV = voidptr

pub const nv_external_compute_queue_spec_version = 1
pub const nv_external_compute_queue_extension_name = c'VK_NV_external_compute_queue'
// ExternalComputeQueueDeviceCreateInfoNV extends VkDeviceCreateInfo
pub type ExternalComputeQueueDeviceCreateInfoNV = C.VkExternalComputeQueueDeviceCreateInfoNV

@[typedef]
pub struct C.VkExternalComputeQueueDeviceCreateInfoNV {
pub mut:
	sType                  StructureType = StructureType.external_compute_queue_device_create_info_nv
	pNext                  voidptr       = unsafe { nil }
	reservedExternalQueues u32
}

pub type ExternalComputeQueueCreateInfoNV = C.VkExternalComputeQueueCreateInfoNV

@[typedef]
pub struct C.VkExternalComputeQueueCreateInfoNV {
pub mut:
	sType          StructureType = StructureType.external_compute_queue_create_info_nv
	pNext          voidptr       = unsafe { nil }
	preferredQueue Queue
}

pub type ExternalComputeQueueDataParamsNV = C.VkExternalComputeQueueDataParamsNV

@[typedef]
pub struct C.VkExternalComputeQueueDataParamsNV {
pub mut:
	sType       StructureType = StructureType.external_compute_queue_data_params_nv
	pNext       voidptr       = unsafe { nil }
	deviceIndex u32
}

// PhysicalDeviceExternalComputeQueuePropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceExternalComputeQueuePropertiesNV = C.VkPhysicalDeviceExternalComputeQueuePropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceExternalComputeQueuePropertiesNV {
pub mut:
	sType             StructureType = StructureType.physical_device_external_compute_queue_properties_nv
	pNext             voidptr       = unsafe { nil }
	externalDataSize  u32
	maxExternalQueues u32
}

@[keep_args_alive]
fn C.vkCreateExternalComputeQueueNV(device Device, p_create_info &ExternalComputeQueueCreateInfoNV, p_allocator &AllocationCallbacks, p_external_queue &ExternalComputeQueueNV) Result

pub type PFN_vkCreateExternalComputeQueueNV = fn (device Device, p_create_info &ExternalComputeQueueCreateInfoNV, p_allocator &AllocationCallbacks, p_external_queue &ExternalComputeQueueNV) Result

@[inline]
pub fn create_external_compute_queue_nv(device Device,
	p_create_info &ExternalComputeQueueCreateInfoNV,
	p_allocator &AllocationCallbacks,
	p_external_queue &ExternalComputeQueueNV) Result {
	return C.vkCreateExternalComputeQueueNV(device, p_create_info, p_allocator, p_external_queue)
}

@[keep_args_alive]
fn C.vkDestroyExternalComputeQueueNV(device Device, external_queue ExternalComputeQueueNV, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyExternalComputeQueueNV = fn (device Device, external_queue ExternalComputeQueueNV, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_external_compute_queue_nv(device Device,
	external_queue ExternalComputeQueueNV,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyExternalComputeQueueNV(device, external_queue, p_allocator)
}

@[keep_args_alive]
fn C.vkGetExternalComputeQueueDataNV(external_queue ExternalComputeQueueNV, mut params ExternalComputeQueueDataParamsNV, p_data voidptr)

pub type PFN_vkGetExternalComputeQueueDataNV = fn (external_queue ExternalComputeQueueNV, mut params ExternalComputeQueueDataParamsNV, p_data voidptr)

@[inline]
pub fn get_external_compute_queue_data_nv(external_queue ExternalComputeQueueNV,
	mut params ExternalComputeQueueDataParamsNV,
	p_data voidptr) {
	C.vkGetExternalComputeQueueDataNV(external_queue, mut params, p_data)
}

pub const nv_command_buffer_inheritance_spec_version = 1
pub const nv_command_buffer_inheritance_extension_name = c'VK_NV_command_buffer_inheritance'
// PhysicalDeviceCommandBufferInheritanceFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCommandBufferInheritanceFeaturesNV = C.VkPhysicalDeviceCommandBufferInheritanceFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceCommandBufferInheritanceFeaturesNV {
pub mut:
	sType                    StructureType = StructureType.physical_device_command_buffer_inheritance_features_nv
	pNext                    voidptr       = unsafe { nil }
	commandBufferInheritance Bool32
}

pub const nv_shader_atomic_float16_vector_spec_version = 1
pub const nv_shader_atomic_float16_vector_extension_name = c'VK_NV_shader_atomic_float16_vector'
// PhysicalDeviceShaderAtomicFloat16VectorFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderAtomicFloat16VectorFeaturesNV = C.VkPhysicalDeviceShaderAtomicFloat16VectorFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceShaderAtomicFloat16VectorFeaturesNV {
pub mut:
	sType                      StructureType = StructureType.physical_device_shader_atomic_float16_vector_features_nv
	pNext                      voidptr       = unsafe { nil }
	shaderFloat16VectorAtomics Bool32
}

pub const ext_shader_replicated_composites_spec_version = 1
pub const ext_shader_replicated_composites_extension_name = c'VK_EXT_shader_replicated_composites'
// PhysicalDeviceShaderReplicatedCompositesFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderReplicatedCompositesFeaturesEXT = C.VkPhysicalDeviceShaderReplicatedCompositesFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderReplicatedCompositesFeaturesEXT {
pub mut:
	sType                      StructureType = StructureType.physical_device_shader_replicated_composites_features_ext
	pNext                      voidptr       = unsafe { nil }
	shaderReplicatedComposites Bool32
}

pub const ext_shader_float8_spec_version = 1
pub const ext_shader_float8_extension_name = c'VK_EXT_shader_float8'
// PhysicalDeviceShaderFloat8FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderFloat8FeaturesEXT = C.VkPhysicalDeviceShaderFloat8FeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderFloat8FeaturesEXT {
pub mut:
	sType                         StructureType = StructureType.physical_device_shader_float8_features_ext
	pNext                         voidptr       = unsafe { nil }
	shaderFloat8                  Bool32
	shaderFloat8CooperativeMatrix Bool32
}

pub const nv_ray_tracing_validation_spec_version = 1
pub const nv_ray_tracing_validation_extension_name = c'VK_NV_ray_tracing_validation'
// PhysicalDeviceRayTracingValidationFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRayTracingValidationFeaturesNV = C.VkPhysicalDeviceRayTracingValidationFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceRayTracingValidationFeaturesNV {
pub mut:
	sType                StructureType = StructureType.physical_device_ray_tracing_validation_features_nv
	pNext                voidptr       = unsafe { nil }
	rayTracingValidation Bool32
}

pub const nv_cluster_acceleration_structure_spec_version = 4
pub const nv_cluster_acceleration_structure_extension_name = c'VK_NV_cluster_acceleration_structure'

pub enum ClusterAccelerationStructureTypeNV as u32 {
	clusters_bottom_level     = 0
	triangle_cluster          = 1
	triangle_cluster_template = 2
	max_enum_nv               = max_int
}

pub enum ClusterAccelerationStructureOpTypeNV as u32 {
	move_objects                    = 0
	build_clusters_bottom_level     = 1
	build_triangle_cluster          = 2
	build_triangle_cluster_template = 3
	instantiate_triangle_cluster    = 4
	get_cluster_template_indices    = 5
	max_enum_nv                     = max_int
}

pub enum ClusterAccelerationStructureOpModeNV as u32 {
	implicit_destinations = 0
	explicit_destinations = 1
	compute_sizes         = 2
	max_enum_nv           = max_int
}

pub enum ClusterAccelerationStructureAddressResolutionFlagBitsNV as u32 {
	none                         = 0
	indirected_dst_implicit_data = u32(0x00000001)
	indirected_scratch_data      = u32(0x00000002)
	indirected_dst_address_array = u32(0x00000004)
	indirected_dst_sizes_array   = u32(0x00000008)
	indirected_src_infos_array   = u32(0x00000010)
	indirected_src_infos_count   = u32(0x00000020)
	max_enum_nv                  = max_int
}
pub type ClusterAccelerationStructureAddressResolutionFlagsNV = u32

pub enum ClusterAccelerationStructureClusterFlagBitsNV as u32 {
	allow_disable_opacity_micromaps = u32(0x00000001)
	max_enum_nv                     = max_int
}
pub type ClusterAccelerationStructureClusterFlagsNV = u32

pub enum ClusterAccelerationStructureGeometryFlagBitsNV as u32 {
	cull_disable                   = u32(0x00000001)
	no_duplicate_anyhit_invocation = u32(0x00000002)
	opaque                         = u32(0x00000004)
	max_enum_nv                    = max_int
}
pub type ClusterAccelerationStructureGeometryFlagsNV = u32

pub enum ClusterAccelerationStructureIndexFormatFlagBitsNV as u32 {
	_8          = u32(0x00000001)
	_16         = u32(0x00000002)
	_32         = u32(0x00000004)
	max_enum_nv = max_int
}
pub type ClusterAccelerationStructureIndexFormatFlagsNV = u32

// PhysicalDeviceClusterAccelerationStructureFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceClusterAccelerationStructureFeaturesNV = C.VkPhysicalDeviceClusterAccelerationStructureFeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceClusterAccelerationStructureFeaturesNV {
pub mut:
	sType                        StructureType = StructureType.physical_device_cluster_acceleration_structure_features_nv
	pNext                        voidptr       = unsafe { nil }
	clusterAccelerationStructure Bool32
}

// PhysicalDeviceClusterAccelerationStructurePropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceClusterAccelerationStructurePropertiesNV = C.VkPhysicalDeviceClusterAccelerationStructurePropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceClusterAccelerationStructurePropertiesNV {
pub mut:
	sType                              StructureType = StructureType.physical_device_cluster_acceleration_structure_properties_nv
	pNext                              voidptr       = unsafe { nil }
	maxVerticesPerCluster              u32
	maxTrianglesPerCluster             u32
	clusterScratchByteAlignment        u32
	clusterByteAlignment               u32
	clusterTemplateByteAlignment       u32
	clusterBottomLevelByteAlignment    u32
	clusterTemplateBoundsByteAlignment u32
	maxClusterGeometryIndex            u32
}

pub type ClusterAccelerationStructureClustersBottomLevelInputNV = C.VkClusterAccelerationStructureClustersBottomLevelInputNV

@[typedef]
pub struct C.VkClusterAccelerationStructureClustersBottomLevelInputNV {
pub mut:
	sType                                   StructureType = StructureType.cluster_acceleration_structure_clusters_bottom_level_input_nv
	pNext                                   voidptr       = unsafe { nil }
	maxTotalClusterCount                    u32
	maxClusterCountPerAccelerationStructure u32
}

pub type ClusterAccelerationStructureTriangleClusterInputNV = C.VkClusterAccelerationStructureTriangleClusterInputNV

@[typedef]
pub struct C.VkClusterAccelerationStructureTriangleClusterInputNV {
pub mut:
	sType                         StructureType = StructureType.cluster_acceleration_structure_triangle_cluster_input_nv
	pNext                         voidptr       = unsafe { nil }
	vertexFormat                  Format
	maxGeometryIndexValue         u32
	maxClusterUniqueGeometryCount u32
	maxClusterTriangleCount       u32
	maxClusterVertexCount         u32
	maxTotalTriangleCount         u32
	maxTotalVertexCount           u32
	minPositionTruncateBitCount   u32
}

pub type ClusterAccelerationStructureMoveObjectsInputNV = C.VkClusterAccelerationStructureMoveObjectsInputNV

@[typedef]
pub struct C.VkClusterAccelerationStructureMoveObjectsInputNV {
pub mut:
	sType         StructureType = StructureType.cluster_acceleration_structure_move_objects_input_nv
	pNext         voidptr       = unsafe { nil }
	type          ClusterAccelerationStructureTypeNV
	noMoveOverlap Bool32
	maxMovedBytes DeviceSize
}

pub type ClusterAccelerationStructureOpInputNV = C.VkClusterAccelerationStructureOpInputNV

@[typedef]
pub union C.VkClusterAccelerationStructureOpInputNV {
pub mut:
	pClustersBottomLevel &ClusterAccelerationStructureClustersBottomLevelInputNV
	pTriangleClusters    &ClusterAccelerationStructureTriangleClusterInputNV
	pMoveObjects         &ClusterAccelerationStructureMoveObjectsInputNV
}

pub type ClusterAccelerationStructureInputInfoNV = C.VkClusterAccelerationStructureInputInfoNV

@[typedef]
pub struct C.VkClusterAccelerationStructureInputInfoNV {
pub mut:
	sType                         StructureType = StructureType.cluster_acceleration_structure_input_info_nv
	pNext                         voidptr       = unsafe { nil }
	maxAccelerationStructureCount u32
	flags                         BuildAccelerationStructureFlagsKHR
	opType                        ClusterAccelerationStructureOpTypeNV
	opMode                        ClusterAccelerationStructureOpModeNV
	opInput                       ClusterAccelerationStructureOpInputNV
}

pub type StridedDeviceAddressRegionKHR = C.VkStridedDeviceAddressRegionKHR

@[typedef]
pub struct C.VkStridedDeviceAddressRegionKHR {
pub mut:
	deviceAddress DeviceAddress
	stride        DeviceSize
	size          DeviceSize
}

pub type ClusterAccelerationStructureCommandsInfoNV = C.VkClusterAccelerationStructureCommandsInfoNV

@[typedef]
pub struct C.VkClusterAccelerationStructureCommandsInfoNV {
pub mut:
	sType                  StructureType = StructureType.cluster_acceleration_structure_commands_info_nv
	pNext                  voidptr       = unsafe { nil }
	input                  ClusterAccelerationStructureInputInfoNV
	dstImplicitData        DeviceAddress
	scratchData            DeviceAddress
	dstAddressesArray      StridedDeviceAddressRegionKHR
	dstSizesArray          StridedDeviceAddressRegionKHR
	srcInfosArray          StridedDeviceAddressRegionKHR
	srcInfosCount          DeviceAddress
	addressResolutionFlags ClusterAccelerationStructureAddressResolutionFlagsNV
}

pub type StridedDeviceAddressNV = C.VkStridedDeviceAddressNV

@[typedef]
pub struct C.VkStridedDeviceAddressNV {
pub mut:
	startAddress  DeviceAddress
	strideInBytes DeviceSize
}

pub type ClusterAccelerationStructureGeometryIndexAndGeometryFlagsNV = C.VkClusterAccelerationStructureGeometryIndexAndGeometryFlagsNV

@[typedef]
pub struct C.VkClusterAccelerationStructureGeometryIndexAndGeometryFlagsNV {
pub mut:
	geometryIndex u32
	reserved      u32
	geometryFlags u32
}

pub type ClusterAccelerationStructureMoveObjectsInfoNV = C.VkClusterAccelerationStructureMoveObjectsInfoNV

@[typedef]
pub struct C.VkClusterAccelerationStructureMoveObjectsInfoNV {
pub mut:
	srcAccelerationStructure DeviceAddress
}

pub type ClusterAccelerationStructureBuildClustersBottomLevelInfoNV = C.VkClusterAccelerationStructureBuildClustersBottomLevelInfoNV

@[typedef]
pub struct C.VkClusterAccelerationStructureBuildClustersBottomLevelInfoNV {
pub mut:
	clusterReferencesCount  u32
	clusterReferencesStride u32
	clusterReferences       DeviceAddress
}

pub type ClusterAccelerationStructureBuildTriangleClusterInfoNV = C.VkClusterAccelerationStructureBuildTriangleClusterInfoNV

@[typedef]
pub struct C.VkClusterAccelerationStructureBuildTriangleClusterInfoNV {
pub mut:
	clusterID                         u32
	clusterFlags                      ClusterAccelerationStructureClusterFlagsNV
	triangleCount                     u32
	vertexCount                       u32
	positionTruncateBitCount          u32
	indexType                         u32
	opacityMicromapIndexType          u32
	baseGeometryIndexAndGeometryFlags ClusterAccelerationStructureGeometryIndexAndGeometryFlagsNV
	indexBufferStride                 u16
	vertexBufferStride                u16
	geometryIndexAndFlagsBufferStride u16
	opacityMicromapIndexBufferStride  u16
	indexBuffer                       DeviceAddress
	vertexBuffer                      DeviceAddress
	geometryIndexAndFlagsBuffer       DeviceAddress
	opacityMicromapArray              DeviceAddress
	opacityMicromapIndexBuffer        DeviceAddress
}

pub type ClusterAccelerationStructureBuildTriangleClusterTemplateInfoNV = C.VkClusterAccelerationStructureBuildTriangleClusterTemplateInfoNV

@[typedef]
pub struct C.VkClusterAccelerationStructureBuildTriangleClusterTemplateInfoNV {
pub mut:
	clusterID                         u32
	clusterFlags                      ClusterAccelerationStructureClusterFlagsNV
	triangleCount                     u32
	vertexCount                       u32
	positionTruncateBitCount          u32
	indexType                         u32
	opacityMicromapIndexType          u32
	baseGeometryIndexAndGeometryFlags ClusterAccelerationStructureGeometryIndexAndGeometryFlagsNV
	indexBufferStride                 u16
	vertexBufferStride                u16
	geometryIndexAndFlagsBufferStride u16
	opacityMicromapIndexBufferStride  u16
	indexBuffer                       DeviceAddress
	vertexBuffer                      DeviceAddress
	geometryIndexAndFlagsBuffer       DeviceAddress
	opacityMicromapArray              DeviceAddress
	opacityMicromapIndexBuffer        DeviceAddress
	instantiationBoundingBoxLimit     DeviceAddress
}

pub type ClusterAccelerationStructureInstantiateClusterInfoNV = C.VkClusterAccelerationStructureInstantiateClusterInfoNV

@[typedef]
pub struct C.VkClusterAccelerationStructureInstantiateClusterInfoNV {
pub mut:
	clusterIdOffset        u32
	geometryIndexOffset    u32
	reserved               u32
	clusterTemplateAddress DeviceAddress
	vertexBuffer           StridedDeviceAddressNV
}

pub type ClusterAccelerationStructureGetTemplateIndicesInfoNV = C.VkClusterAccelerationStructureGetTemplateIndicesInfoNV

@[typedef]
pub struct C.VkClusterAccelerationStructureGetTemplateIndicesInfoNV {
pub mut:
	clusterTemplateAddress DeviceAddress
}

pub type AccelerationStructureBuildSizesInfoKHR = C.VkAccelerationStructureBuildSizesInfoKHR

@[typedef]
pub struct C.VkAccelerationStructureBuildSizesInfoKHR {
pub mut:
	sType                     StructureType = StructureType.acceleration_structure_build_sizes_info_khr
	pNext                     voidptr       = unsafe { nil }
	accelerationStructureSize DeviceSize
	updateScratchSize         DeviceSize
	buildScratchSize          DeviceSize
}

// RayTracingPipelineClusterAccelerationStructureCreateInfoNV extends VkRayTracingPipelineCreateInfoKHR
pub type RayTracingPipelineClusterAccelerationStructureCreateInfoNV = C.VkRayTracingPipelineClusterAccelerationStructureCreateInfoNV

@[typedef]
pub struct C.VkRayTracingPipelineClusterAccelerationStructureCreateInfoNV {
pub mut:
	sType                             StructureType = StructureType.ray_tracing_pipeline_cluster_acceleration_structure_create_info_nv
	pNext                             voidptr       = unsafe { nil }
	allowClusterAccelerationStructure Bool32
}

@[keep_args_alive]
fn C.vkGetClusterAccelerationStructureBuildSizesNV(device Device, p_info &ClusterAccelerationStructureInputInfoNV, mut p_size_info AccelerationStructureBuildSizesInfoKHR)

pub type PFN_vkGetClusterAccelerationStructureBuildSizesNV = fn (device Device, p_info &ClusterAccelerationStructureInputInfoNV, mut p_size_info AccelerationStructureBuildSizesInfoKHR)

@[inline]
pub fn get_cluster_acceleration_structure_build_sizes_nv(device Device,
	p_info &ClusterAccelerationStructureInputInfoNV,
	mut p_size_info AccelerationStructureBuildSizesInfoKHR) {
	C.vkGetClusterAccelerationStructureBuildSizesNV(device, p_info, mut p_size_info)
}

@[keep_args_alive]
fn C.vkCmdBuildClusterAccelerationStructureIndirectNV(command_buffer CommandBuffer, p_command_infos &ClusterAccelerationStructureCommandsInfoNV)

pub type PFN_vkCmdBuildClusterAccelerationStructureIndirectNV = fn (command_buffer CommandBuffer, p_command_infos &ClusterAccelerationStructureCommandsInfoNV)

@[inline]
pub fn cmd_build_cluster_acceleration_structure_indirect_nv(command_buffer CommandBuffer,
	p_command_infos &ClusterAccelerationStructureCommandsInfoNV) {
	C.vkCmdBuildClusterAccelerationStructureIndirectNV(command_buffer, p_command_infos)
}

pub const nv_partitioned_acceleration_structure_spec_version = 1
pub const nv_partitioned_acceleration_structure_extension_name = c'VK_NV_partitioned_acceleration_structure'
pub const partitioned_acceleration_structure_partition_index_global_nv = ~u32(0)

pub enum PartitionedAccelerationStructureOpTypeNV as u32 {
	write_instance              = 0
	update_instance             = 1
	write_partition_translation = 2
	max_enum_nv                 = max_int
}

pub enum PartitionedAccelerationStructureInstanceFlagBitsNV as u32 {
	triangle_facing_cull_disable = u32(0x00000001)
	triangle_flip_facing         = u32(0x00000002)
	force_opaque                 = u32(0x00000004)
	force_no_opaque              = u32(0x00000008)
	enable_explicit_bounding_box = u32(0x00000010)
	max_enum_nv                  = max_int
}
pub type PartitionedAccelerationStructureInstanceFlagsNV = u32

// PhysicalDevicePartitionedAccelerationStructureFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePartitionedAccelerationStructureFeaturesNV = C.VkPhysicalDevicePartitionedAccelerationStructureFeaturesNV

@[typedef]
pub struct C.VkPhysicalDevicePartitionedAccelerationStructureFeaturesNV {
pub mut:
	sType                            StructureType = StructureType.physical_device_partitioned_acceleration_structure_features_nv
	pNext                            voidptr       = unsafe { nil }
	partitionedAccelerationStructure Bool32
}

// PhysicalDevicePartitionedAccelerationStructurePropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDevicePartitionedAccelerationStructurePropertiesNV = C.VkPhysicalDevicePartitionedAccelerationStructurePropertiesNV

@[typedef]
pub struct C.VkPhysicalDevicePartitionedAccelerationStructurePropertiesNV {
pub mut:
	sType             StructureType = StructureType.physical_device_partitioned_acceleration_structure_properties_nv
	pNext             voidptr       = unsafe { nil }
	maxPartitionCount u32
}

// PartitionedAccelerationStructureFlagsNV extends VkPartitionedAccelerationStructureInstancesInputNV
pub type PartitionedAccelerationStructureFlagsNV = C.VkPartitionedAccelerationStructureFlagsNV

@[typedef]
pub struct C.VkPartitionedAccelerationStructureFlagsNV {
pub mut:
	sType                      StructureType = StructureType.partitioned_acceleration_structure_flags_nv
	pNext                      voidptr       = unsafe { nil }
	enablePartitionTranslation Bool32
}

pub type BuildPartitionedAccelerationStructureIndirectCommandNV = C.VkBuildPartitionedAccelerationStructureIndirectCommandNV

@[typedef]
pub struct C.VkBuildPartitionedAccelerationStructureIndirectCommandNV {
pub mut:
	opType   PartitionedAccelerationStructureOpTypeNV
	argCount u32
	argData  StridedDeviceAddressNV
}

pub type PartitionedAccelerationStructureWriteInstanceDataNV = C.VkPartitionedAccelerationStructureWriteInstanceDataNV

@[typedef]
pub struct C.VkPartitionedAccelerationStructureWriteInstanceDataNV {
pub mut:
	transform                           TransformMatrixKHR
	explicitAABB                        [6]f32
	instanceID                          u32
	instanceMask                        u32
	instanceContributionToHitGroupIndex u32
	instanceFlags                       PartitionedAccelerationStructureInstanceFlagsNV
	instanceIndex                       u32
	partitionIndex                      u32
	accelerationStructure               DeviceAddress
}

pub type PartitionedAccelerationStructureUpdateInstanceDataNV = C.VkPartitionedAccelerationStructureUpdateInstanceDataNV

@[typedef]
pub struct C.VkPartitionedAccelerationStructureUpdateInstanceDataNV {
pub mut:
	instanceIndex                       u32
	instanceContributionToHitGroupIndex u32
	accelerationStructure               DeviceAddress
}

pub type PartitionedAccelerationStructureWritePartitionTranslationDataNV = C.VkPartitionedAccelerationStructureWritePartitionTranslationDataNV

@[typedef]
pub struct C.VkPartitionedAccelerationStructureWritePartitionTranslationDataNV {
pub mut:
	partitionIndex       u32
	partitionTranslation [3]f32
}

// WriteDescriptorSetPartitionedAccelerationStructureNV extends VkWriteDescriptorSet
pub type WriteDescriptorSetPartitionedAccelerationStructureNV = C.VkWriteDescriptorSetPartitionedAccelerationStructureNV

@[typedef]
pub struct C.VkWriteDescriptorSetPartitionedAccelerationStructureNV {
pub mut:
	sType                      StructureType = StructureType.write_descriptor_set_partitioned_acceleration_structure_nv
	pNext                      voidptr       = unsafe { nil }
	accelerationStructureCount u32
	pAccelerationStructures    &DeviceAddress
}

pub type PartitionedAccelerationStructureInstancesInputNV = C.VkPartitionedAccelerationStructureInstancesInputNV

@[typedef]
pub struct C.VkPartitionedAccelerationStructureInstancesInputNV {
pub mut:
	sType                             StructureType = StructureType.partitioned_acceleration_structure_instances_input_nv
	pNext                             voidptr       = unsafe { nil }
	flags                             BuildAccelerationStructureFlagsKHR
	instanceCount                     u32
	maxInstancePerPartitionCount      u32
	partitionCount                    u32
	maxInstanceInGlobalPartitionCount u32
}

pub type BuildPartitionedAccelerationStructureInfoNV = C.VkBuildPartitionedAccelerationStructureInfoNV

@[typedef]
pub struct C.VkBuildPartitionedAccelerationStructureInfoNV {
pub mut:
	sType                        StructureType = StructureType.build_partitioned_acceleration_structure_info_nv
	pNext                        voidptr       = unsafe { nil }
	input                        PartitionedAccelerationStructureInstancesInputNV
	srcAccelerationStructureData DeviceAddress
	dstAccelerationStructureData DeviceAddress
	scratchData                  DeviceAddress
	srcInfos                     DeviceAddress
	srcInfosCount                DeviceAddress
}

@[keep_args_alive]
fn C.vkGetPartitionedAccelerationStructuresBuildSizesNV(device Device, p_info &PartitionedAccelerationStructureInstancesInputNV, mut p_size_info AccelerationStructureBuildSizesInfoKHR)

pub type PFN_vkGetPartitionedAccelerationStructuresBuildSizesNV = fn (device Device, p_info &PartitionedAccelerationStructureInstancesInputNV, mut p_size_info AccelerationStructureBuildSizesInfoKHR)

@[inline]
pub fn get_partitioned_acceleration_structures_build_sizes_nv(device Device,
	p_info &PartitionedAccelerationStructureInstancesInputNV,
	mut p_size_info AccelerationStructureBuildSizesInfoKHR) {
	C.vkGetPartitionedAccelerationStructuresBuildSizesNV(device, p_info, mut p_size_info)
}

@[keep_args_alive]
fn C.vkCmdBuildPartitionedAccelerationStructuresNV(command_buffer CommandBuffer, p_build_info &BuildPartitionedAccelerationStructureInfoNV)

pub type PFN_vkCmdBuildPartitionedAccelerationStructuresNV = fn (command_buffer CommandBuffer, p_build_info &BuildPartitionedAccelerationStructureInfoNV)

@[inline]
pub fn cmd_build_partitioned_acceleration_structures_nv(command_buffer CommandBuffer,
	p_build_info &BuildPartitionedAccelerationStructureInfoNV) {
	C.vkCmdBuildPartitionedAccelerationStructuresNV(command_buffer, p_build_info)
}

// Pointer to VkIndirectExecutionSetEXT_T
pub type IndirectExecutionSetEXT = voidptr

// Pointer to VkIndirectCommandsLayoutEXT_T
pub type IndirectCommandsLayoutEXT = voidptr

pub const ext_device_generated_commands_spec_version = 1
pub const ext_device_generated_commands_extension_name = c'VK_EXT_device_generated_commands'

pub enum IndirectExecutionSetInfoTypeEXT as u32 {
	pipelines      = 0
	shader_objects = 1
	max_enum_ext   = max_int
}

pub enum IndirectCommandsTokenTypeEXT as u32 {
	execution_set            = 0
	push_constant            = 1
	sequence_index           = 2
	index_buffer             = 3
	vertex_buffer            = 4
	draw_indexed             = 5
	draw                     = 6
	draw_indexed_count       = 7
	draw_count               = 8
	dispatch                 = 9
	draw_mesh_tasks_nv       = 1000202002
	draw_mesh_tasks_count_nv = 1000202003
	draw_mesh_tasks          = 1000328000
	draw_mesh_tasks_count    = 1000328001
	trace_rays2              = 1000386004
	max_enum_ext             = max_int
}

pub enum IndirectCommandsInputModeFlagBitsEXT as u32 {
	vulkan_index_buffer = u32(0x00000001)
	dxgi_index_buffer   = u32(0x00000002)
	max_enum_ext        = max_int
}
pub type IndirectCommandsInputModeFlagsEXT = u32

pub enum IndirectCommandsLayoutUsageFlagBitsEXT as u32 {
	explicit_preprocess = u32(0x00000001)
	unordered_sequences = u32(0x00000002)
	max_enum_ext        = max_int
}
pub type IndirectCommandsLayoutUsageFlagsEXT = u32

// PhysicalDeviceDeviceGeneratedCommandsFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDeviceGeneratedCommandsFeaturesEXT = C.VkPhysicalDeviceDeviceGeneratedCommandsFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDeviceGeneratedCommandsFeaturesEXT {
pub mut:
	sType                          StructureType = StructureType.physical_device_device_generated_commands_features_ext
	pNext                          voidptr       = unsafe { nil }
	deviceGeneratedCommands        Bool32
	dynamicGeneratedPipelineLayout Bool32
}

// PhysicalDeviceDeviceGeneratedCommandsPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceDeviceGeneratedCommandsPropertiesEXT = C.VkPhysicalDeviceDeviceGeneratedCommandsPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDeviceGeneratedCommandsPropertiesEXT {
pub mut:
	sType                                                StructureType = StructureType.physical_device_device_generated_commands_properties_ext
	pNext                                                voidptr       = unsafe { nil }
	maxIndirectPipelineCount                             u32
	maxIndirectShaderObjectCount                         u32
	maxIndirectSequenceCount                             u32
	maxIndirectCommandsTokenCount                        u32
	maxIndirectCommandsTokenOffset                       u32
	maxIndirectCommandsIndirectStride                    u32
	supportedIndirectCommandsInputModes                  IndirectCommandsInputModeFlagsEXT
	supportedIndirectCommandsShaderStages                ShaderStageFlags
	supportedIndirectCommandsShaderStagesPipelineBinding ShaderStageFlags
	supportedIndirectCommandsShaderStagesShaderBinding   ShaderStageFlags
	deviceGeneratedCommandsTransformFeedback             Bool32
	deviceGeneratedCommandsMultiDrawIndirectCount        Bool32
}

pub type GeneratedCommandsMemoryRequirementsInfoEXT = C.VkGeneratedCommandsMemoryRequirementsInfoEXT

@[typedef]
pub struct C.VkGeneratedCommandsMemoryRequirementsInfoEXT {
pub mut:
	sType                  StructureType = StructureType.generated_commands_memory_requirements_info_ext
	pNext                  voidptr       = unsafe { nil }
	indirectExecutionSet   IndirectExecutionSetEXT
	indirectCommandsLayout IndirectCommandsLayoutEXT
	maxSequenceCount       u32
	maxDrawCount           u32
}

pub type IndirectExecutionSetPipelineInfoEXT = C.VkIndirectExecutionSetPipelineInfoEXT

@[typedef]
pub struct C.VkIndirectExecutionSetPipelineInfoEXT {
pub mut:
	sType            StructureType = StructureType.indirect_execution_set_pipeline_info_ext
	pNext            voidptr       = unsafe { nil }
	initialPipeline  Pipeline
	maxPipelineCount u32
}

pub type IndirectExecutionSetShaderLayoutInfoEXT = C.VkIndirectExecutionSetShaderLayoutInfoEXT

@[typedef]
pub struct C.VkIndirectExecutionSetShaderLayoutInfoEXT {
pub mut:
	sType          StructureType = StructureType.indirect_execution_set_shader_layout_info_ext
	pNext          voidptr       = unsafe { nil }
	setLayoutCount u32
	pSetLayouts    &DescriptorSetLayout
}

pub type IndirectExecutionSetShaderInfoEXT = C.VkIndirectExecutionSetShaderInfoEXT

@[typedef]
pub struct C.VkIndirectExecutionSetShaderInfoEXT {
pub mut:
	sType                  StructureType = StructureType.indirect_execution_set_shader_info_ext
	pNext                  voidptr       = unsafe { nil }
	shaderCount            u32
	pInitialShaders        &ShaderEXT
	pSetLayoutInfos        &IndirectExecutionSetShaderLayoutInfoEXT
	maxShaderCount         u32
	pushConstantRangeCount u32
	pPushConstantRanges    &PushConstantRange
}

pub type IndirectExecutionSetInfoEXT = C.VkIndirectExecutionSetInfoEXT

@[typedef]
pub union C.VkIndirectExecutionSetInfoEXT {
pub mut:
	pPipelineInfo &IndirectExecutionSetPipelineInfoEXT
	pShaderInfo   &IndirectExecutionSetShaderInfoEXT
}

pub type IndirectExecutionSetCreateInfoEXT = C.VkIndirectExecutionSetCreateInfoEXT

@[typedef]
pub struct C.VkIndirectExecutionSetCreateInfoEXT {
pub mut:
	sType StructureType = StructureType.indirect_execution_set_create_info_ext
	pNext voidptr       = unsafe { nil }
	type  IndirectExecutionSetInfoTypeEXT
	info  IndirectExecutionSetInfoEXT
}

pub type GeneratedCommandsInfoEXT = C.VkGeneratedCommandsInfoEXT

@[typedef]
pub struct C.VkGeneratedCommandsInfoEXT {
pub mut:
	sType                  StructureType = StructureType.generated_commands_info_ext
	pNext                  voidptr       = unsafe { nil }
	shaderStages           ShaderStageFlags
	indirectExecutionSet   IndirectExecutionSetEXT
	indirectCommandsLayout IndirectCommandsLayoutEXT
	indirectAddress        DeviceAddress
	indirectAddressSize    DeviceSize
	preprocessAddress      DeviceAddress
	preprocessSize         DeviceSize
	maxSequenceCount       u32
	sequenceCountAddress   DeviceAddress
	maxDrawCount           u32
}

pub type WriteIndirectExecutionSetPipelineEXT = C.VkWriteIndirectExecutionSetPipelineEXT

@[typedef]
pub struct C.VkWriteIndirectExecutionSetPipelineEXT {
pub mut:
	sType    StructureType = StructureType.write_indirect_execution_set_pipeline_ext
	pNext    voidptr       = unsafe { nil }
	index    u32
	pipeline Pipeline
}

pub type IndirectCommandsPushConstantTokenEXT = C.VkIndirectCommandsPushConstantTokenEXT

@[typedef]
pub struct C.VkIndirectCommandsPushConstantTokenEXT {
pub mut:
	updateRange PushConstantRange
}

pub type IndirectCommandsVertexBufferTokenEXT = C.VkIndirectCommandsVertexBufferTokenEXT

@[typedef]
pub struct C.VkIndirectCommandsVertexBufferTokenEXT {
pub mut:
	vertexBindingUnit u32
}

pub type IndirectCommandsIndexBufferTokenEXT = C.VkIndirectCommandsIndexBufferTokenEXT

@[typedef]
pub struct C.VkIndirectCommandsIndexBufferTokenEXT {
pub mut:
	mode IndirectCommandsInputModeFlagBitsEXT
}

pub type IndirectCommandsExecutionSetTokenEXT = C.VkIndirectCommandsExecutionSetTokenEXT

@[typedef]
pub struct C.VkIndirectCommandsExecutionSetTokenEXT {
pub mut:
	type         IndirectExecutionSetInfoTypeEXT
	shaderStages ShaderStageFlags
}

pub type IndirectCommandsTokenDataEXT = C.VkIndirectCommandsTokenDataEXT

@[typedef]
pub union C.VkIndirectCommandsTokenDataEXT {
pub mut:
	pPushConstant &IndirectCommandsPushConstantTokenEXT
	pVertexBuffer &IndirectCommandsVertexBufferTokenEXT
	pIndexBuffer  &IndirectCommandsIndexBufferTokenEXT
	pExecutionSet &IndirectCommandsExecutionSetTokenEXT
}

pub type IndirectCommandsLayoutTokenEXT = C.VkIndirectCommandsLayoutTokenEXT

@[typedef]
pub struct C.VkIndirectCommandsLayoutTokenEXT {
pub mut:
	sType  StructureType = StructureType.indirect_commands_layout_token_ext
	pNext  voidptr       = unsafe { nil }
	type   IndirectCommandsTokenTypeEXT
	data   IndirectCommandsTokenDataEXT
	offset u32
}

pub type IndirectCommandsLayoutCreateInfoEXT = C.VkIndirectCommandsLayoutCreateInfoEXT

@[typedef]
pub struct C.VkIndirectCommandsLayoutCreateInfoEXT {
pub mut:
	sType          StructureType = StructureType.indirect_commands_layout_create_info_ext
	pNext          voidptr       = unsafe { nil }
	flags          IndirectCommandsLayoutUsageFlagsEXT
	shaderStages   ShaderStageFlags
	indirectStride u32
	pipelineLayout PipelineLayout
	tokenCount     u32
	pTokens        &IndirectCommandsLayoutTokenEXT
}

pub type DrawIndirectCountIndirectCommandEXT = C.VkDrawIndirectCountIndirectCommandEXT

@[typedef]
pub struct C.VkDrawIndirectCountIndirectCommandEXT {
pub mut:
	bufferAddress DeviceAddress
	stride        u32
	commandCount  u32
}

pub type BindVertexBufferIndirectCommandEXT = C.VkBindVertexBufferIndirectCommandEXT

@[typedef]
pub struct C.VkBindVertexBufferIndirectCommandEXT {
pub mut:
	bufferAddress DeviceAddress
	size          u32
	stride        u32
}

pub type BindIndexBufferIndirectCommandEXT = C.VkBindIndexBufferIndirectCommandEXT

@[typedef]
pub struct C.VkBindIndexBufferIndirectCommandEXT {
pub mut:
	bufferAddress DeviceAddress
	size          u32
	indexType     IndexType
}

// GeneratedCommandsPipelineInfoEXT extends VkGeneratedCommandsInfoEXT,VkGeneratedCommandsMemoryRequirementsInfoEXT
pub type GeneratedCommandsPipelineInfoEXT = C.VkGeneratedCommandsPipelineInfoEXT

@[typedef]
pub struct C.VkGeneratedCommandsPipelineInfoEXT {
pub mut:
	sType    StructureType = StructureType.generated_commands_pipeline_info_ext
	pNext    voidptr       = unsafe { nil }
	pipeline Pipeline
}

// GeneratedCommandsShaderInfoEXT extends VkGeneratedCommandsInfoEXT,VkGeneratedCommandsMemoryRequirementsInfoEXT
pub type GeneratedCommandsShaderInfoEXT = C.VkGeneratedCommandsShaderInfoEXT

@[typedef]
pub struct C.VkGeneratedCommandsShaderInfoEXT {
pub mut:
	sType       StructureType = StructureType.generated_commands_shader_info_ext
	pNext       voidptr       = unsafe { nil }
	shaderCount u32
	pShaders    &ShaderEXT
}

pub type WriteIndirectExecutionSetShaderEXT = C.VkWriteIndirectExecutionSetShaderEXT

@[typedef]
pub struct C.VkWriteIndirectExecutionSetShaderEXT {
pub mut:
	sType  StructureType = StructureType.write_indirect_execution_set_shader_ext
	pNext  voidptr       = unsafe { nil }
	index  u32
	shader ShaderEXT
}

@[keep_args_alive]
fn C.vkGetGeneratedCommandsMemoryRequirementsEXT(device Device, p_info &GeneratedCommandsMemoryRequirementsInfoEXT, mut p_memory_requirements MemoryRequirements2)

pub type PFN_vkGetGeneratedCommandsMemoryRequirementsEXT = fn (device Device, p_info &GeneratedCommandsMemoryRequirementsInfoEXT, mut p_memory_requirements MemoryRequirements2)

@[inline]
pub fn get_generated_commands_memory_requirements_ext(device Device,
	p_info &GeneratedCommandsMemoryRequirementsInfoEXT,
	mut p_memory_requirements MemoryRequirements2) {
	C.vkGetGeneratedCommandsMemoryRequirementsEXT(device, p_info, mut p_memory_requirements)
}

@[keep_args_alive]
fn C.vkCmdPreprocessGeneratedCommandsEXT(command_buffer CommandBuffer, p_generated_commands_info &GeneratedCommandsInfoEXT, state_command_buffer CommandBuffer)

pub type PFN_vkCmdPreprocessGeneratedCommandsEXT = fn (command_buffer CommandBuffer, p_generated_commands_info &GeneratedCommandsInfoEXT, state_command_buffer CommandBuffer)

@[inline]
pub fn cmd_preprocess_generated_commands_ext(command_buffer CommandBuffer,
	p_generated_commands_info &GeneratedCommandsInfoEXT,
	state_command_buffer CommandBuffer) {
	C.vkCmdPreprocessGeneratedCommandsEXT(command_buffer, p_generated_commands_info, state_command_buffer)
}

@[keep_args_alive]
fn C.vkCmdExecuteGeneratedCommandsEXT(command_buffer CommandBuffer, is_preprocessed Bool32, p_generated_commands_info &GeneratedCommandsInfoEXT)

pub type PFN_vkCmdExecuteGeneratedCommandsEXT = fn (command_buffer CommandBuffer, is_preprocessed Bool32, p_generated_commands_info &GeneratedCommandsInfoEXT)

@[inline]
pub fn cmd_execute_generated_commands_ext(command_buffer CommandBuffer,
	is_preprocessed Bool32,
	p_generated_commands_info &GeneratedCommandsInfoEXT) {
	C.vkCmdExecuteGeneratedCommandsEXT(command_buffer, is_preprocessed, p_generated_commands_info)
}

@[keep_args_alive]
fn C.vkCreateIndirectCommandsLayoutEXT(device Device, p_create_info &IndirectCommandsLayoutCreateInfoEXT, p_allocator &AllocationCallbacks, p_indirect_commands_layout &IndirectCommandsLayoutEXT) Result

pub type PFN_vkCreateIndirectCommandsLayoutEXT = fn (device Device, p_create_info &IndirectCommandsLayoutCreateInfoEXT, p_allocator &AllocationCallbacks, p_indirect_commands_layout &IndirectCommandsLayoutEXT) Result

@[inline]
pub fn create_indirect_commands_layout_ext(device Device,
	p_create_info &IndirectCommandsLayoutCreateInfoEXT,
	p_allocator &AllocationCallbacks,
	p_indirect_commands_layout &IndirectCommandsLayoutEXT) Result {
	return C.vkCreateIndirectCommandsLayoutEXT(device, p_create_info, p_allocator, p_indirect_commands_layout)
}

@[keep_args_alive]
fn C.vkDestroyIndirectCommandsLayoutEXT(device Device, indirect_commands_layout IndirectCommandsLayoutEXT, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyIndirectCommandsLayoutEXT = fn (device Device, indirect_commands_layout IndirectCommandsLayoutEXT, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_indirect_commands_layout_ext(device Device,
	indirect_commands_layout IndirectCommandsLayoutEXT,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyIndirectCommandsLayoutEXT(device, indirect_commands_layout, p_allocator)
}

@[keep_args_alive]
fn C.vkCreateIndirectExecutionSetEXT(device Device, p_create_info &IndirectExecutionSetCreateInfoEXT, p_allocator &AllocationCallbacks, p_indirect_execution_set &IndirectExecutionSetEXT) Result

pub type PFN_vkCreateIndirectExecutionSetEXT = fn (device Device, p_create_info &IndirectExecutionSetCreateInfoEXT, p_allocator &AllocationCallbacks, p_indirect_execution_set &IndirectExecutionSetEXT) Result

@[inline]
pub fn create_indirect_execution_set_ext(device Device,
	p_create_info &IndirectExecutionSetCreateInfoEXT,
	p_allocator &AllocationCallbacks,
	p_indirect_execution_set &IndirectExecutionSetEXT) Result {
	return C.vkCreateIndirectExecutionSetEXT(device, p_create_info, p_allocator, p_indirect_execution_set)
}

@[keep_args_alive]
fn C.vkDestroyIndirectExecutionSetEXT(device Device, indirect_execution_set IndirectExecutionSetEXT, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyIndirectExecutionSetEXT = fn (device Device, indirect_execution_set IndirectExecutionSetEXT, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_indirect_execution_set_ext(device Device,
	indirect_execution_set IndirectExecutionSetEXT,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyIndirectExecutionSetEXT(device, indirect_execution_set, p_allocator)
}

@[keep_args_alive]
fn C.vkUpdateIndirectExecutionSetPipelineEXT(device Device, indirect_execution_set IndirectExecutionSetEXT, execution_set_write_count u32, p_execution_set_writes &WriteIndirectExecutionSetPipelineEXT)

pub type PFN_vkUpdateIndirectExecutionSetPipelineEXT = fn (device Device, indirect_execution_set IndirectExecutionSetEXT, execution_set_write_count u32, p_execution_set_writes &WriteIndirectExecutionSetPipelineEXT)

@[inline]
pub fn update_indirect_execution_set_pipeline_ext(device Device,
	indirect_execution_set IndirectExecutionSetEXT,
	execution_set_write_count u32,
	p_execution_set_writes &WriteIndirectExecutionSetPipelineEXT) {
	C.vkUpdateIndirectExecutionSetPipelineEXT(device, indirect_execution_set, execution_set_write_count,
		p_execution_set_writes)
}

@[keep_args_alive]
fn C.vkUpdateIndirectExecutionSetShaderEXT(device Device, indirect_execution_set IndirectExecutionSetEXT, execution_set_write_count u32, p_execution_set_writes &WriteIndirectExecutionSetShaderEXT)

pub type PFN_vkUpdateIndirectExecutionSetShaderEXT = fn (device Device, indirect_execution_set IndirectExecutionSetEXT, execution_set_write_count u32, p_execution_set_writes &WriteIndirectExecutionSetShaderEXT)

@[inline]
pub fn update_indirect_execution_set_shader_ext(device Device,
	indirect_execution_set IndirectExecutionSetEXT,
	execution_set_write_count u32,
	p_execution_set_writes &WriteIndirectExecutionSetShaderEXT) {
	C.vkUpdateIndirectExecutionSetShaderEXT(device, indirect_execution_set, execution_set_write_count,
		p_execution_set_writes)
}

pub const mesa_image_alignment_control_spec_version = 1
pub const mesa_image_alignment_control_extension_name = c'VK_MESA_image_alignment_control'
// PhysicalDeviceImageAlignmentControlFeaturesMESA extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceImageAlignmentControlFeaturesMESA = C.VkPhysicalDeviceImageAlignmentControlFeaturesMESA

@[typedef]
pub struct C.VkPhysicalDeviceImageAlignmentControlFeaturesMESA {
pub mut:
	sType                 StructureType = StructureType.physical_device_image_alignment_control_features_mesa
	pNext                 voidptr       = unsafe { nil }
	imageAlignmentControl Bool32
}

// PhysicalDeviceImageAlignmentControlPropertiesMESA extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceImageAlignmentControlPropertiesMESA = C.VkPhysicalDeviceImageAlignmentControlPropertiesMESA

@[typedef]
pub struct C.VkPhysicalDeviceImageAlignmentControlPropertiesMESA {
pub mut:
	sType                       StructureType = StructureType.physical_device_image_alignment_control_properties_mesa
	pNext                       voidptr       = unsafe { nil }
	supportedImageAlignmentMask u32
}

// ImageAlignmentControlCreateInfoMESA extends VkImageCreateInfo
pub type ImageAlignmentControlCreateInfoMESA = C.VkImageAlignmentControlCreateInfoMESA

@[typedef]
pub struct C.VkImageAlignmentControlCreateInfoMESA {
pub mut:
	sType                     StructureType = StructureType.image_alignment_control_create_info_mesa
	pNext                     voidptr       = unsafe { nil }
	maximumRequestedAlignment u32
}

pub const ext_depth_clamp_control_spec_version = 1
pub const ext_depth_clamp_control_extension_name = c'VK_EXT_depth_clamp_control'
// PhysicalDeviceDepthClampControlFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceDepthClampControlFeaturesEXT = C.VkPhysicalDeviceDepthClampControlFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceDepthClampControlFeaturesEXT {
pub mut:
	sType             StructureType = StructureType.physical_device_depth_clamp_control_features_ext
	pNext             voidptr       = unsafe { nil }
	depthClampControl Bool32
}

// PipelineViewportDepthClampControlCreateInfoEXT extends VkPipelineViewportStateCreateInfo
pub type PipelineViewportDepthClampControlCreateInfoEXT = C.VkPipelineViewportDepthClampControlCreateInfoEXT

@[typedef]
pub struct C.VkPipelineViewportDepthClampControlCreateInfoEXT {
pub mut:
	sType            StructureType = StructureType.pipeline_viewport_depth_clamp_control_create_info_ext
	pNext            voidptr       = unsafe { nil }
	depthClampMode   DepthClampModeEXT
	pDepthClampRange &DepthClampRangeEXT
}

pub type OHNativeWindow = C.OHNativeWindow

@[typedef]
pub struct C.OHNativeWindow {}

pub const ohos_surface_spec_version = 1
pub const ohos_surface_extension_name = c'VK_OHOS_surface'

pub type SurfaceCreateFlagsOHOS = u32
pub type SurfaceCreateInfoOHOS = C.VkSurfaceCreateInfoOHOS

@[typedef]
pub struct C.VkSurfaceCreateInfoOHOS {
pub mut:
	sType  StructureType = StructureType.surface_create_info_ohos
	pNext  voidptr       = unsafe { nil }
	flags  SurfaceCreateFlagsOHOS
	window &OHNativeWindow
}

@[keep_args_alive]
fn C.vkCreateSurfaceOHOS(instance Instance, p_create_info &SurfaceCreateInfoOHOS, p_allocator &AllocationCallbacks, p_surface &SurfaceKHR) Result

pub type PFN_vkCreateSurfaceOHOS = fn (instance Instance, p_create_info &SurfaceCreateInfoOHOS, p_allocator &AllocationCallbacks, p_surface &SurfaceKHR) Result

@[inline]
pub fn create_surface_ohos(instance Instance,
	p_create_info &SurfaceCreateInfoOHOS,
	p_allocator &AllocationCallbacks,
	p_surface &SurfaceKHR) Result {
	return C.vkCreateSurfaceOHOS(instance, p_create_info, p_allocator, p_surface)
}

pub type OHBufferHandle = C.OHBufferHandle

@[typedef]
pub struct C.OHBufferHandle {}

pub const ohos_native_buffer_spec_version = 1
pub const ohos_native_buffer_extension_name = c'VK_OHOS_native_buffer'

pub enum SwapchainImageUsageFlagBitsOHOS as u32 {
	shared        = u32(0x00000001)
	max_enum_ohos = max_int
}
pub type SwapchainImageUsageFlagsOHOS = u32

// NativeBufferOHOS extends VkImageCreateInfo,VkBindImageMemoryInfo
pub type NativeBufferOHOS = C.VkNativeBufferOHOS

@[typedef]
pub struct C.VkNativeBufferOHOS {
pub mut:
	sType  StructureType = StructureType.native_buffer_ohos
	pNext  voidptr       = unsafe { nil }
	handle &OHBufferHandle
}

// SwapchainImageCreateInfoOHOS extends VkImageCreateInfo
pub type SwapchainImageCreateInfoOHOS = C.VkSwapchainImageCreateInfoOHOS

@[typedef]
pub struct C.VkSwapchainImageCreateInfoOHOS {
pub mut:
	sType StructureType = StructureType.swapchain_image_create_info_ohos
	pNext voidptr       = unsafe { nil }
	usage SwapchainImageUsageFlagsOHOS
}

// PhysicalDevicePresentationPropertiesOHOS extends VkPhysicalDeviceProperties2
pub type PhysicalDevicePresentationPropertiesOHOS = C.VkPhysicalDevicePresentationPropertiesOHOS

@[typedef]
pub struct C.VkPhysicalDevicePresentationPropertiesOHOS {
pub mut:
	sType       StructureType = StructureType.physical_device_presentation_properties_ohos
	pNext       voidptr       = unsafe { nil }
	sharedImage Bool32
}

@[keep_args_alive]
fn C.vkGetSwapchainGrallocUsageOHOS(device Device, format Format, image_usage ImageUsageFlags, gralloc_usage &u64) Result

pub type PFN_vkGetSwapchainGrallocUsageOHOS = fn (device Device, format Format, image_usage ImageUsageFlags, gralloc_usage &u64) Result

@[inline]
pub fn get_swapchain_gralloc_usage_ohos(device Device,
	format Format,
	image_usage ImageUsageFlags,
	gralloc_usage &u64) Result {
	return C.vkGetSwapchainGrallocUsageOHOS(device, format, image_usage, gralloc_usage)
}

@[keep_args_alive]
fn C.vkAcquireImageOHOS(device Device, image Image, native_fence_fd i32, semaphore Semaphore, fence Fence) Result

pub type PFN_vkAcquireImageOHOS = fn (device Device, image Image, native_fence_fd i32, semaphore Semaphore, fence Fence) Result

@[inline]
pub fn acquire_image_ohos(device Device,
	image Image,
	native_fence_fd i32,
	semaphore Semaphore,
	fence Fence) Result {
	return C.vkAcquireImageOHOS(device, image, native_fence_fd, semaphore, fence)
}

@[keep_args_alive]
fn C.vkQueueSignalReleaseImageOHOS(queue Queue, wait_semaphore_count u32, p_wait_semaphores &Semaphore, image Image, p_native_fence_fd &i32) Result

pub type PFN_vkQueueSignalReleaseImageOHOS = fn (queue Queue, wait_semaphore_count u32, p_wait_semaphores &Semaphore, image Image, p_native_fence_fd &i32) Result

@[inline]
pub fn queue_signal_release_image_ohos(queue Queue,
	wait_semaphore_count u32,
	p_wait_semaphores &Semaphore,
	image Image,
	p_native_fence_fd &i32) Result {
	return C.vkQueueSignalReleaseImageOHOS(queue, wait_semaphore_count, p_wait_semaphores,
		image, p_native_fence_fd)
}

pub const huawei_hdr_vivid_spec_version = 1
pub const huawei_hdr_vivid_extension_name = c'VK_HAWEI_hdr_vivid'
// PhysicalDeviceHdrVividFeaturesHUAWEI extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceHdrVividFeaturesHUAWEI = C.VkPhysicalDeviceHdrVividFeaturesHUAWEI

@[typedef]
pub struct C.VkPhysicalDeviceHdrVividFeaturesHUAWEI {
pub mut:
	sType    StructureType = StructureType.physical_device_hdr_vivid_features_huawei
	pNext    voidptr       = unsafe { nil }
	hdrVivid Bool32
}

// HdrVividDynamicMetadataHUAWEI extends VkHdrMetadataEXT
pub type HdrVividDynamicMetadataHUAWEI = C.VkHdrVividDynamicMetadataHUAWEI

@[typedef]
pub struct C.VkHdrVividDynamicMetadataHUAWEI {
pub mut:
	sType               StructureType = StructureType.hdr_vivid_dynamic_metadata_huawei
	pNext               voidptr       = unsafe { nil }
	dynamicMetadataSize usize
	pDynamicMetadata    voidptr
}

pub const nv_cooperative_matrix_2_spec_version = 1
pub const nv_cooperative_matrix_2_extension_name = c'VK_NV_cooperative_matrix2'

pub type CooperativeMatrixFlexibleDimensionsPropertiesNV = C.VkCooperativeMatrixFlexibleDimensionsPropertiesNV

@[typedef]
pub struct C.VkCooperativeMatrixFlexibleDimensionsPropertiesNV {
pub mut:
	sType                  StructureType = StructureType.cooperative_matrix_flexible_dimensions_properties_nv
	pNext                  voidptr       = unsafe { nil }
	MGranularity           u32
	NGranularity           u32
	KGranularity           u32
	AType                  ComponentTypeKHR
	BType                  ComponentTypeKHR
	CType                  ComponentTypeKHR
	ResultType             ComponentTypeKHR
	saturatingAccumulation Bool32
	scope                  ScopeKHR
	workgroupInvocations   u32
}

// PhysicalDeviceCooperativeMatrix2FeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceCooperativeMatrix2FeaturesNV = C.VkPhysicalDeviceCooperativeMatrix2FeaturesNV

@[typedef]
pub struct C.VkPhysicalDeviceCooperativeMatrix2FeaturesNV {
pub mut:
	sType                                 StructureType = StructureType.physical_device_cooperative_matrix2_features_nv
	pNext                                 voidptr       = unsafe { nil }
	cooperativeMatrixWorkgroupScope       Bool32
	cooperativeMatrixFlexibleDimensions   Bool32
	cooperativeMatrixReductions           Bool32
	cooperativeMatrixConversions          Bool32
	cooperativeMatrixPerElementOperations Bool32
	cooperativeMatrixTensorAddressing     Bool32
	cooperativeMatrixBlockLoads           Bool32
}

// PhysicalDeviceCooperativeMatrix2PropertiesNV extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceCooperativeMatrix2PropertiesNV = C.VkPhysicalDeviceCooperativeMatrix2PropertiesNV

@[typedef]
pub struct C.VkPhysicalDeviceCooperativeMatrix2PropertiesNV {
pub mut:
	sType                                               StructureType = StructureType.physical_device_cooperative_matrix2_properties_nv
	pNext                                               voidptr       = unsafe { nil }
	cooperativeMatrixWorkgroupScopeMaxWorkgroupSize     u32
	cooperativeMatrixFlexibleDimensionsMaxDimension     u32
	cooperativeMatrixWorkgroupScopeReservedSharedMemory u32
}

@[keep_args_alive]
fn C.vkGetPhysicalDeviceCooperativeMatrixFlexibleDimensionsPropertiesNV(physical_device PhysicalDevice, p_property_count &u32, mut p_properties CooperativeMatrixFlexibleDimensionsPropertiesNV) Result

pub type PFN_vkGetPhysicalDeviceCooperativeMatrixFlexibleDimensionsPropertiesNV = fn (physical_device PhysicalDevice, p_property_count &u32, mut p_properties CooperativeMatrixFlexibleDimensionsPropertiesNV) Result

@[inline]
pub fn get_physical_device_cooperative_matrix_flexible_dimensions_properties_nv(physical_device PhysicalDevice,
	p_property_count &u32,
	mut p_properties CooperativeMatrixFlexibleDimensionsPropertiesNV) Result {
	return C.vkGetPhysicalDeviceCooperativeMatrixFlexibleDimensionsPropertiesNV(physical_device,
		p_property_count, mut p_properties)
}

pub const arm_pipeline_opacity_micromap_spec_version = 1
pub const arm_pipeline_opacity_micromap_extension_name = c'VK_ARM_pipeline_opacity_micromap'
// PhysicalDevicePipelineOpacityMicromapFeaturesARM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePipelineOpacityMicromapFeaturesARM = C.VkPhysicalDevicePipelineOpacityMicromapFeaturesARM

@[typedef]
pub struct C.VkPhysicalDevicePipelineOpacityMicromapFeaturesARM {
pub mut:
	sType                   StructureType = StructureType.physical_device_pipeline_opacity_micromap_features_arm
	pNext                   voidptr       = unsafe { nil }
	pipelineOpacityMicromap Bool32
}

pub const ext_external_memory_metal_spec_version = 1
pub const ext_external_memory_metal_extension_name = c'VK_EXT_external_memory_metal'
// ImportMemoryMetalHandleInfoEXT extends VkMemoryAllocateInfo
pub type ImportMemoryMetalHandleInfoEXT = C.VkImportMemoryMetalHandleInfoEXT

@[typedef]
pub struct C.VkImportMemoryMetalHandleInfoEXT {
pub mut:
	sType      StructureType = StructureType.import_memory_metal_handle_info_ext
	pNext      voidptr       = unsafe { nil }
	handleType ExternalMemoryHandleTypeFlagBits
	handle     voidptr
}

pub type MemoryMetalHandlePropertiesEXT = C.VkMemoryMetalHandlePropertiesEXT

@[typedef]
pub struct C.VkMemoryMetalHandlePropertiesEXT {
pub mut:
	sType          StructureType = StructureType.memory_metal_handle_properties_ext
	pNext          voidptr       = unsafe { nil }
	memoryTypeBits u32
}

pub type MemoryGetMetalHandleInfoEXT = C.VkMemoryGetMetalHandleInfoEXT

@[typedef]
pub struct C.VkMemoryGetMetalHandleInfoEXT {
pub mut:
	sType      StructureType = StructureType.memory_get_metal_handle_info_ext
	pNext      voidptr       = unsafe { nil }
	memory     DeviceMemory
	handleType ExternalMemoryHandleTypeFlagBits
}

@[keep_args_alive]
fn C.vkGetMemoryMetalHandleEXT(device Device, p_get_metal_handle_info &MemoryGetMetalHandleInfoEXT, p_handle &voidptr) Result

pub type PFN_vkGetMemoryMetalHandleEXT = fn (device Device, p_get_metal_handle_info &MemoryGetMetalHandleInfoEXT, p_handle &voidptr) Result

@[inline]
pub fn get_memory_metal_handle_ext(device Device,
	p_get_metal_handle_info &MemoryGetMetalHandleInfoEXT,
	p_handle &voidptr) Result {
	return C.vkGetMemoryMetalHandleEXT(device, p_get_metal_handle_info, p_handle)
}

@[keep_args_alive]
fn C.vkGetMemoryMetalHandlePropertiesEXT(device Device, handle_type ExternalMemoryHandleTypeFlagBits, p_handle voidptr, mut p_memory_metal_handle_properties MemoryMetalHandlePropertiesEXT) Result

pub type PFN_vkGetMemoryMetalHandlePropertiesEXT = fn (device Device, handle_type ExternalMemoryHandleTypeFlagBits, p_handle voidptr, mut p_memory_metal_handle_properties MemoryMetalHandlePropertiesEXT) Result

@[inline]
pub fn get_memory_metal_handle_properties_ext(device Device,
	handle_type ExternalMemoryHandleTypeFlagBits,
	p_handle voidptr,
	mut p_memory_metal_handle_properties MemoryMetalHandlePropertiesEXT) Result {
	return C.vkGetMemoryMetalHandlePropertiesEXT(device, handle_type, p_handle, mut p_memory_metal_handle_properties)
}

pub const ext_vertex_attribute_robustness_spec_version = 1
pub const ext_vertex_attribute_robustness_extension_name = c'VK_EXT_vertex_attribute_robustness'
// PhysicalDeviceVertexAttributeRobustnessFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceVertexAttributeRobustnessFeaturesEXT = C.VkPhysicalDeviceVertexAttributeRobustnessFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceVertexAttributeRobustnessFeaturesEXT {
pub mut:
	sType                     StructureType = StructureType.physical_device_vertex_attribute_robustness_features_ext
	pNext                     voidptr       = unsafe { nil }
	vertexAttributeRobustness Bool32
}

pub const arm_format_pack_spec_version = 1
pub const arm_format_pack_extension_name = c'VK_ARM_format_pack'
// PhysicalDeviceFormatPackFeaturesARM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceFormatPackFeaturesARM = C.VkPhysicalDeviceFormatPackFeaturesARM

@[typedef]
pub struct C.VkPhysicalDeviceFormatPackFeaturesARM {
pub mut:
	sType      StructureType = StructureType.physical_device_format_pack_features_arm
	pNext      voidptr       = unsafe { nil }
	formatPack Bool32
}

pub const valve_fragment_density_map_layered_spec_version = 1
pub const valve_fragment_density_map_layered_extension_name = c'VK_VAVE_fragment_density_map_layered'
// PhysicalDeviceFragmentDensityMapLayeredFeaturesVALVE extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceFragmentDensityMapLayeredFeaturesVALVE = C.VkPhysicalDeviceFragmentDensityMapLayeredFeaturesVALVE

@[typedef]
pub struct C.VkPhysicalDeviceFragmentDensityMapLayeredFeaturesVALVE {
pub mut:
	sType                     StructureType = StructureType.physical_device_fragment_density_map_layered_features_valve
	pNext                     voidptr       = unsafe { nil }
	fragmentDensityMapLayered Bool32
}

// PhysicalDeviceFragmentDensityMapLayeredPropertiesVALVE extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceFragmentDensityMapLayeredPropertiesVALVE = C.VkPhysicalDeviceFragmentDensityMapLayeredPropertiesVALVE

@[typedef]
pub struct C.VkPhysicalDeviceFragmentDensityMapLayeredPropertiesVALVE {
pub mut:
	sType                       StructureType = StructureType.physical_device_fragment_density_map_layered_properties_valve
	pNext                       voidptr       = unsafe { nil }
	maxFragmentDensityMapLayers u32
}

// PipelineFragmentDensityMapLayeredCreateInfoVALVE extends VkGraphicsPipelineCreateInfo
pub type PipelineFragmentDensityMapLayeredCreateInfoVALVE = C.VkPipelineFragmentDensityMapLayeredCreateInfoVALVE

@[typedef]
pub struct C.VkPipelineFragmentDensityMapLayeredCreateInfoVALVE {
pub mut:
	sType                       StructureType = StructureType.pipeline_fragment_density_map_layered_create_info_valve
	pNext                       voidptr       = unsafe { nil }
	maxFragmentDensityMapLayers u32
}

pub const nv_present_metering_spec_version = 1
pub const nv_present_metering_extension_name = c'VK_NV_present_metering'
// SetPresentConfigNV extends VkPresentInfoKHR
pub type SetPresentConfigNV = C.VkSetPresentConfigNV

@[typedef]
pub struct C.VkSetPresentConfigNV {
pub mut:
	sType                 StructureType
	pNext                 voidptr = unsafe { nil }
	numFramesPerBatch     u32
	presentConfigFeedback u32
}

// PhysicalDevicePresentMeteringFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePresentMeteringFeaturesNV = C.VkPhysicalDevicePresentMeteringFeaturesNV

@[typedef]
pub struct C.VkPhysicalDevicePresentMeteringFeaturesNV {
pub mut:
	sType           StructureType
	pNext           voidptr = unsafe { nil }
	presentMetering Bool32
}

pub const ext_fragment_density_map_offset_spec_version = 1
pub const ext_fragment_density_map_offset_extension_name = c'VK_EXT_fragment_density_map_offset'

pub type RenderingEndInfoEXT = C.VkRenderingEndInfoKHR

@[keep_args_alive]
fn C.vkCmdEndRendering2EXT(command_buffer CommandBuffer, p_rendering_end_info &RenderingEndInfoKHR)

pub type PFN_vkCmdEndRendering2EXT = fn (command_buffer CommandBuffer, p_rendering_end_info &RenderingEndInfoKHR)

@[inline]
pub fn cmd_end_rendering2_ext(command_buffer CommandBuffer,
	p_rendering_end_info &RenderingEndInfoKHR) {
	C.vkCmdEndRendering2EXT(command_buffer, p_rendering_end_info)
}

pub const ext_zero_initialize_device_memory_spec_version = 1
pub const ext_zero_initialize_device_memory_extension_name = c'VK_EXT_zero_initialize_device_memory'
// PhysicalDeviceZeroInitializeDeviceMemoryFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceZeroInitializeDeviceMemoryFeaturesEXT = C.VkPhysicalDeviceZeroInitializeDeviceMemoryFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceZeroInitializeDeviceMemoryFeaturesEXT {
pub mut:
	sType                      StructureType = StructureType.physical_device_zero_initialize_device_memory_features_ext
	pNext                      voidptr       = unsafe { nil }
	zeroInitializeDeviceMemory Bool32
}

pub const ext_shader_64bit_indexing_spec_version = 1
pub const ext_shader_64bit_indexing_extension_name = c'VK_EXT_shader_64bit_indexing'
// PhysicalDeviceShader64BitIndexingFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShader64BitIndexingFeaturesEXT = C.VkPhysicalDeviceShader64BitIndexingFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShader64BitIndexingFeaturesEXT {
pub mut:
	sType               StructureType = StructureType.physical_device_shader64_bit_indexing_features_ext
	pNext               voidptr       = unsafe { nil }
	shader64BitIndexing Bool32
}

pub const sec_pipeline_cache_incremental_mode_spec_version = 1
pub const sec_pipeline_cache_incremental_mode_extension_name = c'VK_SEC_pipeline_cache_incremental_mode'
// PhysicalDevicePipelineCacheIncrementalModeFeaturesSEC extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDevicePipelineCacheIncrementalModeFeaturesSEC = C.VkPhysicalDevicePipelineCacheIncrementalModeFeaturesSEC

@[typedef]
pub struct C.VkPhysicalDevicePipelineCacheIncrementalModeFeaturesSEC {
pub mut:
	sType                        StructureType = StructureType.physical_device_pipeline_cache_incremental_mode_features_sec
	pNext                        voidptr       = unsafe { nil }
	pipelineCacheIncrementalMode Bool32
}

pub const ext_shader_uniform_buffer_unsized_array_spec_version = 1
pub const ext_shader_uniform_buffer_unsized_array_extension_name = c'VK_EXT_shader_uniform_buffer_unsized_array'
// PhysicalDeviceShaderUniformBufferUnsizedArrayFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceShaderUniformBufferUnsizedArrayFeaturesEXT = C.VkPhysicalDeviceShaderUniformBufferUnsizedArrayFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceShaderUniformBufferUnsizedArrayFeaturesEXT {
pub mut:
	sType                           StructureType = StructureType.physical_device_shader_uniform_buffer_unsized_array_features_ext
	pNext                           voidptr       = unsafe { nil }
	shaderUniformBufferUnsizedArray Bool32
}

pub const khr_acceleration_structure_spec_version = 13
pub const khr_acceleration_structure_extension_name = c'VK_KHR_acceleration_structure'

pub enum BuildAccelerationStructureModeKHR as u32 {
	build        = 0
	update       = 1
	max_enum_khr = max_int
}

pub enum AccelerationStructureCreateFlagBitsKHR as u32 {
	device_address_capture_replay            = u32(0x00000001)
	descriptor_buffer_capture_replay_bit_ext = u32(0x00000008)
	motion_bit_nv                            = u32(0x00000004)
	max_enum_khr                             = max_int
}
pub type AccelerationStructureCreateFlagsKHR = u32
pub type AccelerationStructureBuildRangeInfoKHR = C.VkAccelerationStructureBuildRangeInfoKHR

@[typedef]
pub struct C.VkAccelerationStructureBuildRangeInfoKHR {
pub mut:
	primitiveCount  u32
	primitiveOffset u32
	firstVertex     u32
	transformOffset u32
}

pub type AccelerationStructureGeometryTrianglesDataKHR = C.VkAccelerationStructureGeometryTrianglesDataKHR

@[typedef]
pub struct C.VkAccelerationStructureGeometryTrianglesDataKHR {
pub mut:
	sType         StructureType = StructureType.acceleration_structure_geometry_triangles_data_khr
	pNext         voidptr       = unsafe { nil }
	vertexFormat  Format
	vertexData    DeviceOrHostAddressConstKHR
	vertexStride  DeviceSize
	maxVertex     u32
	indexType     IndexType
	indexData     DeviceOrHostAddressConstKHR
	transformData DeviceOrHostAddressConstKHR
}

pub type AccelerationStructureGeometryAabbsDataKHR = C.VkAccelerationStructureGeometryAabbsDataKHR

@[typedef]
pub struct C.VkAccelerationStructureGeometryAabbsDataKHR {
pub mut:
	sType  StructureType = StructureType.acceleration_structure_geometry_aabbs_data_khr
	pNext  voidptr       = unsafe { nil }
	data   DeviceOrHostAddressConstKHR
	stride DeviceSize
}

pub type AccelerationStructureGeometryInstancesDataKHR = C.VkAccelerationStructureGeometryInstancesDataKHR

@[typedef]
pub struct C.VkAccelerationStructureGeometryInstancesDataKHR {
pub mut:
	sType           StructureType = StructureType.acceleration_structure_geometry_instances_data_khr
	pNext           voidptr       = unsafe { nil }
	arrayOfPointers Bool32
	data            DeviceOrHostAddressConstKHR
}

pub type AccelerationStructureGeometryDataKHR = C.VkAccelerationStructureGeometryDataKHR

@[typedef]
pub union C.VkAccelerationStructureGeometryDataKHR {
pub mut:
	triangles AccelerationStructureGeometryTrianglesDataKHR
	aabbs     AccelerationStructureGeometryAabbsDataKHR
	instances AccelerationStructureGeometryInstancesDataKHR
}

pub type AccelerationStructureGeometryKHR = C.VkAccelerationStructureGeometryKHR

@[typedef]
pub struct C.VkAccelerationStructureGeometryKHR {
pub mut:
	sType        StructureType = StructureType.acceleration_structure_geometry_khr
	pNext        voidptr       = unsafe { nil }
	geometryType GeometryTypeKHR
	geometry     AccelerationStructureGeometryDataKHR
	flags        GeometryFlagsKHR
}

pub type AccelerationStructureBuildGeometryInfoKHR = C.VkAccelerationStructureBuildGeometryInfoKHR

@[typedef]
pub struct C.VkAccelerationStructureBuildGeometryInfoKHR {
pub mut:
	sType                    StructureType = StructureType.acceleration_structure_build_geometry_info_khr
	pNext                    voidptr       = unsafe { nil }
	type                     AccelerationStructureTypeKHR
	flags                    BuildAccelerationStructureFlagsKHR
	mode                     BuildAccelerationStructureModeKHR
	srcAccelerationStructure AccelerationStructureKHR
	dstAccelerationStructure AccelerationStructureKHR
	geometryCount            u32
	pGeometries              &AccelerationStructureGeometryKHR
	ppGeometries             &&AccelerationStructureGeometryKHR
	scratchData              DeviceOrHostAddressKHR
}

pub type AccelerationStructureCreateInfoKHR = C.VkAccelerationStructureCreateInfoKHR

@[typedef]
pub struct C.VkAccelerationStructureCreateInfoKHR {
pub mut:
	sType         StructureType = StructureType.acceleration_structure_create_info_khr
	pNext         voidptr       = unsafe { nil }
	createFlags   AccelerationStructureCreateFlagsKHR
	buffer        Buffer
	offset        DeviceSize
	size          DeviceSize
	type          AccelerationStructureTypeKHR
	deviceAddress DeviceAddress
}

// WriteDescriptorSetAccelerationStructureKHR extends VkWriteDescriptorSet
pub type WriteDescriptorSetAccelerationStructureKHR = C.VkWriteDescriptorSetAccelerationStructureKHR

@[typedef]
pub struct C.VkWriteDescriptorSetAccelerationStructureKHR {
pub mut:
	sType                      StructureType = StructureType.write_descriptor_set_acceleration_structure_khr
	pNext                      voidptr       = unsafe { nil }
	accelerationStructureCount u32
	pAccelerationStructures    &AccelerationStructureKHR
}

// PhysicalDeviceAccelerationStructureFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceAccelerationStructureFeaturesKHR = C.VkPhysicalDeviceAccelerationStructureFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceAccelerationStructureFeaturesKHR {
pub mut:
	sType                                                 StructureType = StructureType.physical_device_acceleration_structure_features_khr
	pNext                                                 voidptr       = unsafe { nil }
	accelerationStructure                                 Bool32
	accelerationStructureCaptureReplay                    Bool32
	accelerationStructureIndirectBuild                    Bool32
	accelerationStructureHostCommands                     Bool32
	descriptorBindingAccelerationStructureUpdateAfterBind Bool32
}

// PhysicalDeviceAccelerationStructurePropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceAccelerationStructurePropertiesKHR = C.VkPhysicalDeviceAccelerationStructurePropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceAccelerationStructurePropertiesKHR {
pub mut:
	sType                                                      StructureType = StructureType.physical_device_acceleration_structure_properties_khr
	pNext                                                      voidptr       = unsafe { nil }
	maxGeometryCount                                           u64
	maxInstanceCount                                           u64
	maxPrimitiveCount                                          u64
	maxPerStageDescriptorAccelerationStructures                u32
	maxPerStageDescriptorUpdateAfterBindAccelerationStructures u32
	maxDescriptorSetAccelerationStructures                     u32
	maxDescriptorSetUpdateAfterBindAccelerationStructures      u32
	minAccelerationStructureScratchOffsetAlignment             u32
}

pub type AccelerationStructureDeviceAddressInfoKHR = C.VkAccelerationStructureDeviceAddressInfoKHR

@[typedef]
pub struct C.VkAccelerationStructureDeviceAddressInfoKHR {
pub mut:
	sType                 StructureType = StructureType.acceleration_structure_device_address_info_khr
	pNext                 voidptr       = unsafe { nil }
	accelerationStructure AccelerationStructureKHR
}

pub type AccelerationStructureVersionInfoKHR = C.VkAccelerationStructureVersionInfoKHR

@[typedef]
pub struct C.VkAccelerationStructureVersionInfoKHR {
pub mut:
	sType        StructureType = StructureType.acceleration_structure_version_info_khr
	pNext        voidptr       = unsafe { nil }
	pVersionData &u8
}

pub type CopyAccelerationStructureToMemoryInfoKHR = C.VkCopyAccelerationStructureToMemoryInfoKHR

@[typedef]
pub struct C.VkCopyAccelerationStructureToMemoryInfoKHR {
pub mut:
	sType StructureType = StructureType.copy_acceleration_structure_to_memory_info_khr
	pNext voidptr       = unsafe { nil }
	src   AccelerationStructureKHR
	dst   DeviceOrHostAddressKHR
	mode  CopyAccelerationStructureModeKHR
}

pub type CopyMemoryToAccelerationStructureInfoKHR = C.VkCopyMemoryToAccelerationStructureInfoKHR

@[typedef]
pub struct C.VkCopyMemoryToAccelerationStructureInfoKHR {
pub mut:
	sType StructureType = StructureType.copy_memory_to_acceleration_structure_info_khr
	pNext voidptr       = unsafe { nil }
	src   DeviceOrHostAddressConstKHR
	dst   AccelerationStructureKHR
	mode  CopyAccelerationStructureModeKHR
}

pub type CopyAccelerationStructureInfoKHR = C.VkCopyAccelerationStructureInfoKHR

@[typedef]
pub struct C.VkCopyAccelerationStructureInfoKHR {
pub mut:
	sType StructureType = StructureType.copy_acceleration_structure_info_khr
	pNext voidptr       = unsafe { nil }
	src   AccelerationStructureKHR
	dst   AccelerationStructureKHR
	mode  CopyAccelerationStructureModeKHR
}

@[keep_args_alive]
fn C.vkCreateAccelerationStructureKHR(device Device, p_create_info &AccelerationStructureCreateInfoKHR, p_allocator &AllocationCallbacks, p_acceleration_structure &AccelerationStructureKHR) Result

pub type PFN_vkCreateAccelerationStructureKHR = fn (device Device, p_create_info &AccelerationStructureCreateInfoKHR, p_allocator &AllocationCallbacks, p_acceleration_structure &AccelerationStructureKHR) Result

@[inline]
pub fn create_acceleration_structure_khr(device Device,
	p_create_info &AccelerationStructureCreateInfoKHR,
	p_allocator &AllocationCallbacks,
	p_acceleration_structure &AccelerationStructureKHR) Result {
	return C.vkCreateAccelerationStructureKHR(device, p_create_info, p_allocator, p_acceleration_structure)
}

@[keep_args_alive]
fn C.vkDestroyAccelerationStructureKHR(device Device, acceleration_structure AccelerationStructureKHR, p_allocator &AllocationCallbacks)

pub type PFN_vkDestroyAccelerationStructureKHR = fn (device Device, acceleration_structure AccelerationStructureKHR, p_allocator &AllocationCallbacks)

@[inline]
pub fn destroy_acceleration_structure_khr(device Device,
	acceleration_structure AccelerationStructureKHR,
	p_allocator &AllocationCallbacks) {
	C.vkDestroyAccelerationStructureKHR(device, acceleration_structure, p_allocator)
}

@[keep_args_alive]
fn C.vkCmdBuildAccelerationStructuresKHR(command_buffer CommandBuffer, info_count u32, p_infos &AccelerationStructureBuildGeometryInfoKHR, pp_build_range_infos &&AccelerationStructureBuildRangeInfoKHR)

pub type PFN_vkCmdBuildAccelerationStructuresKHR = fn (command_buffer CommandBuffer, info_count u32, p_infos &AccelerationStructureBuildGeometryInfoKHR, pp_build_range_infos &&AccelerationStructureBuildRangeInfoKHR)

@[inline]
pub fn cmd_build_acceleration_structures_khr(command_buffer CommandBuffer,
	info_count u32,
	p_infos &AccelerationStructureBuildGeometryInfoKHR,
	pp_build_range_infos &&AccelerationStructureBuildRangeInfoKHR) {
	C.vkCmdBuildAccelerationStructuresKHR(command_buffer, info_count, p_infos, pp_build_range_infos)
}

@[keep_args_alive]
fn C.vkCmdBuildAccelerationStructuresIndirectKHR(command_buffer CommandBuffer, info_count u32, p_infos &AccelerationStructureBuildGeometryInfoKHR, p_indirect_device_addresses &DeviceAddress, p_indirect_strides &u32, pp_max_primitive_counts &&u32)

pub type PFN_vkCmdBuildAccelerationStructuresIndirectKHR = fn (command_buffer CommandBuffer, info_count u32, p_infos &AccelerationStructureBuildGeometryInfoKHR, p_indirect_device_addresses &DeviceAddress, p_indirect_strides &u32, pp_max_primitive_counts &&u32)

@[inline]
pub fn cmd_build_acceleration_structures_indirect_khr(command_buffer CommandBuffer,
	info_count u32,
	p_infos &AccelerationStructureBuildGeometryInfoKHR,
	p_indirect_device_addresses &DeviceAddress,
	p_indirect_strides &u32,
	pp_max_primitive_counts &&u32) {
	C.vkCmdBuildAccelerationStructuresIndirectKHR(command_buffer, info_count, p_infos,
		p_indirect_device_addresses, p_indirect_strides, pp_max_primitive_counts)
}

@[keep_args_alive]
fn C.vkBuildAccelerationStructuresKHR(device Device, deferred_operation DeferredOperationKHR, info_count u32, p_infos &AccelerationStructureBuildGeometryInfoKHR, pp_build_range_infos &&AccelerationStructureBuildRangeInfoKHR) Result

pub type PFN_vkBuildAccelerationStructuresKHR = fn (device Device, deferred_operation DeferredOperationKHR, info_count u32, p_infos &AccelerationStructureBuildGeometryInfoKHR, pp_build_range_infos &&AccelerationStructureBuildRangeInfoKHR) Result

@[inline]
pub fn build_acceleration_structures_khr(device Device,
	deferred_operation DeferredOperationKHR,
	info_count u32,
	p_infos &AccelerationStructureBuildGeometryInfoKHR,
	pp_build_range_infos &&AccelerationStructureBuildRangeInfoKHR) Result {
	return C.vkBuildAccelerationStructuresKHR(device, deferred_operation, info_count,
		p_infos, pp_build_range_infos)
}

@[keep_args_alive]
fn C.vkCopyAccelerationStructureKHR(device Device, deferred_operation DeferredOperationKHR, p_info &CopyAccelerationStructureInfoKHR) Result

pub type PFN_vkCopyAccelerationStructureKHR = fn (device Device, deferred_operation DeferredOperationKHR, p_info &CopyAccelerationStructureInfoKHR) Result

@[inline]
pub fn copy_acceleration_structure_khr(device Device,
	deferred_operation DeferredOperationKHR,
	p_info &CopyAccelerationStructureInfoKHR) Result {
	return C.vkCopyAccelerationStructureKHR(device, deferred_operation, p_info)
}

@[keep_args_alive]
fn C.vkCopyAccelerationStructureToMemoryKHR(device Device, deferred_operation DeferredOperationKHR, p_info &CopyAccelerationStructureToMemoryInfoKHR) Result

pub type PFN_vkCopyAccelerationStructureToMemoryKHR = fn (device Device, deferred_operation DeferredOperationKHR, p_info &CopyAccelerationStructureToMemoryInfoKHR) Result

@[inline]
pub fn copy_acceleration_structure_to_memory_khr(device Device,
	deferred_operation DeferredOperationKHR,
	p_info &CopyAccelerationStructureToMemoryInfoKHR) Result {
	return C.vkCopyAccelerationStructureToMemoryKHR(device, deferred_operation, p_info)
}

@[keep_args_alive]
fn C.vkCopyMemoryToAccelerationStructureKHR(device Device, deferred_operation DeferredOperationKHR, p_info &CopyMemoryToAccelerationStructureInfoKHR) Result

pub type PFN_vkCopyMemoryToAccelerationStructureKHR = fn (device Device, deferred_operation DeferredOperationKHR, p_info &CopyMemoryToAccelerationStructureInfoKHR) Result

@[inline]
pub fn copy_memory_to_acceleration_structure_khr(device Device,
	deferred_operation DeferredOperationKHR,
	p_info &CopyMemoryToAccelerationStructureInfoKHR) Result {
	return C.vkCopyMemoryToAccelerationStructureKHR(device, deferred_operation, p_info)
}

@[keep_args_alive]
fn C.vkWriteAccelerationStructuresPropertiesKHR(device Device, acceleration_structure_count u32, p_acceleration_structures &AccelerationStructureKHR, query_type QueryType, data_size usize, p_data voidptr, stride usize) Result

pub type PFN_vkWriteAccelerationStructuresPropertiesKHR = fn (device Device, acceleration_structure_count u32, p_acceleration_structures &AccelerationStructureKHR, query_type QueryType, data_size usize, p_data voidptr, stride usize) Result

@[inline]
pub fn write_acceleration_structures_properties_khr(device Device,
	acceleration_structure_count u32,
	p_acceleration_structures &AccelerationStructureKHR,
	query_type QueryType,
	data_size usize,
	p_data voidptr,
	stride usize) Result {
	return C.vkWriteAccelerationStructuresPropertiesKHR(device, acceleration_structure_count,
		p_acceleration_structures, query_type, data_size, p_data, stride)
}

@[keep_args_alive]
fn C.vkCmdCopyAccelerationStructureKHR(command_buffer CommandBuffer, p_info &CopyAccelerationStructureInfoKHR)

pub type PFN_vkCmdCopyAccelerationStructureKHR = fn (command_buffer CommandBuffer, p_info &CopyAccelerationStructureInfoKHR)

@[inline]
pub fn cmd_copy_acceleration_structure_khr(command_buffer CommandBuffer,
	p_info &CopyAccelerationStructureInfoKHR) {
	C.vkCmdCopyAccelerationStructureKHR(command_buffer, p_info)
}

@[keep_args_alive]
fn C.vkCmdCopyAccelerationStructureToMemoryKHR(command_buffer CommandBuffer, p_info &CopyAccelerationStructureToMemoryInfoKHR)

pub type PFN_vkCmdCopyAccelerationStructureToMemoryKHR = fn (command_buffer CommandBuffer, p_info &CopyAccelerationStructureToMemoryInfoKHR)

@[inline]
pub fn cmd_copy_acceleration_structure_to_memory_khr(command_buffer CommandBuffer,
	p_info &CopyAccelerationStructureToMemoryInfoKHR) {
	C.vkCmdCopyAccelerationStructureToMemoryKHR(command_buffer, p_info)
}

@[keep_args_alive]
fn C.vkCmdCopyMemoryToAccelerationStructureKHR(command_buffer CommandBuffer, p_info &CopyMemoryToAccelerationStructureInfoKHR)

pub type PFN_vkCmdCopyMemoryToAccelerationStructureKHR = fn (command_buffer CommandBuffer, p_info &CopyMemoryToAccelerationStructureInfoKHR)

@[inline]
pub fn cmd_copy_memory_to_acceleration_structure_khr(command_buffer CommandBuffer,
	p_info &CopyMemoryToAccelerationStructureInfoKHR) {
	C.vkCmdCopyMemoryToAccelerationStructureKHR(command_buffer, p_info)
}

@[keep_args_alive]
fn C.vkGetAccelerationStructureDeviceAddressKHR(device Device, p_info &AccelerationStructureDeviceAddressInfoKHR) DeviceAddress

pub type PFN_vkGetAccelerationStructureDeviceAddressKHR = fn (device Device, p_info &AccelerationStructureDeviceAddressInfoKHR) DeviceAddress

@[inline]
pub fn get_acceleration_structure_device_address_khr(device Device,
	p_info &AccelerationStructureDeviceAddressInfoKHR) DeviceAddress {
	return C.vkGetAccelerationStructureDeviceAddressKHR(device, p_info)
}

@[keep_args_alive]
fn C.vkCmdWriteAccelerationStructuresPropertiesKHR(command_buffer CommandBuffer, acceleration_structure_count u32, p_acceleration_structures &AccelerationStructureKHR, query_type QueryType, query_pool QueryPool, first_query u32)

pub type PFN_vkCmdWriteAccelerationStructuresPropertiesKHR = fn (command_buffer CommandBuffer, acceleration_structure_count u32, p_acceleration_structures &AccelerationStructureKHR, query_type QueryType, query_pool QueryPool, first_query u32)

@[inline]
pub fn cmd_write_acceleration_structures_properties_khr(command_buffer CommandBuffer,
	acceleration_structure_count u32,
	p_acceleration_structures &AccelerationStructureKHR,
	query_type QueryType,
	query_pool QueryPool,
	first_query u32) {
	C.vkCmdWriteAccelerationStructuresPropertiesKHR(command_buffer, acceleration_structure_count,
		p_acceleration_structures, query_type, query_pool, first_query)
}

@[keep_args_alive]
fn C.vkGetDeviceAccelerationStructureCompatibilityKHR(device Device, p_version_info &AccelerationStructureVersionInfoKHR, p_compatibility &AccelerationStructureCompatibilityKHR)

pub type PFN_vkGetDeviceAccelerationStructureCompatibilityKHR = fn (device Device, p_version_info &AccelerationStructureVersionInfoKHR, p_compatibility &AccelerationStructureCompatibilityKHR)

@[inline]
pub fn get_device_acceleration_structure_compatibility_khr(device Device,
	p_version_info &AccelerationStructureVersionInfoKHR,
	p_compatibility &AccelerationStructureCompatibilityKHR) {
	C.vkGetDeviceAccelerationStructureCompatibilityKHR(device, p_version_info, p_compatibility)
}

@[keep_args_alive]
fn C.vkGetAccelerationStructureBuildSizesKHR(device Device, build_type AccelerationStructureBuildTypeKHR, p_build_info &AccelerationStructureBuildGeometryInfoKHR, p_max_primitive_counts &u32, mut p_size_info AccelerationStructureBuildSizesInfoKHR)

pub type PFN_vkGetAccelerationStructureBuildSizesKHR = fn (device Device, build_type AccelerationStructureBuildTypeKHR, p_build_info &AccelerationStructureBuildGeometryInfoKHR, p_max_primitive_counts &u32, mut p_size_info AccelerationStructureBuildSizesInfoKHR)

@[inline]
pub fn get_acceleration_structure_build_sizes_khr(device Device,
	build_type AccelerationStructureBuildTypeKHR,
	p_build_info &AccelerationStructureBuildGeometryInfoKHR,
	p_max_primitive_counts &u32,
	mut p_size_info AccelerationStructureBuildSizesInfoKHR) {
	C.vkGetAccelerationStructureBuildSizesKHR(device, build_type, p_build_info, p_max_primitive_counts, mut
		p_size_info)
}

pub const khr_ray_tracing_pipeline_spec_version = 1
pub const khr_ray_tracing_pipeline_extension_name = c'VK_KHR_ray_tracing_pipeline'

pub enum ShaderGroupShaderKHR as u32 {
	general      = 0
	closest_hit  = 1
	any_hit      = 2
	intersection = 3
	max_enum_khr = max_int
}
pub type RayTracingShaderGroupCreateInfoKHR = C.VkRayTracingShaderGroupCreateInfoKHR

@[typedef]
pub struct C.VkRayTracingShaderGroupCreateInfoKHR {
pub mut:
	sType                           StructureType = StructureType.ray_tracing_shader_group_create_info_khr
	pNext                           voidptr       = unsafe { nil }
	type                            RayTracingShaderGroupTypeKHR
	generalShader                   u32
	closestHitShader                u32
	anyHitShader                    u32
	intersectionShader              u32
	pShaderGroupCaptureReplayHandle voidptr
}

pub type RayTracingPipelineInterfaceCreateInfoKHR = C.VkRayTracingPipelineInterfaceCreateInfoKHR

@[typedef]
pub struct C.VkRayTracingPipelineInterfaceCreateInfoKHR {
pub mut:
	sType                          StructureType = StructureType.ray_tracing_pipeline_interface_create_info_khr
	pNext                          voidptr       = unsafe { nil }
	maxPipelineRayPayloadSize      u32
	maxPipelineRayHitAttributeSize u32
}

pub type RayTracingPipelineCreateInfoKHR = C.VkRayTracingPipelineCreateInfoKHR

@[typedef]
pub struct C.VkRayTracingPipelineCreateInfoKHR {
pub mut:
	sType                        StructureType = StructureType.ray_tracing_pipeline_create_info_khr
	pNext                        voidptr       = unsafe { nil }
	flags                        PipelineCreateFlags
	stageCount                   u32
	pStages                      &PipelineShaderStageCreateInfo
	groupCount                   u32
	pGroups                      &RayTracingShaderGroupCreateInfoKHR
	maxPipelineRayRecursionDepth u32
	pLibraryInfo                 &PipelineLibraryCreateInfoKHR
	pLibraryInterface            &RayTracingPipelineInterfaceCreateInfoKHR
	pDynamicState                &PipelineDynamicStateCreateInfo
	layout                       PipelineLayout
	basePipelineHandle           Pipeline
	basePipelineIndex            i32
}

// PhysicalDeviceRayTracingPipelineFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRayTracingPipelineFeaturesKHR = C.VkPhysicalDeviceRayTracingPipelineFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceRayTracingPipelineFeaturesKHR {
pub mut:
	sType                                                 StructureType = StructureType.physical_device_ray_tracing_pipeline_features_khr
	pNext                                                 voidptr       = unsafe { nil }
	rayTracingPipeline                                    Bool32
	rayTracingPipelineShaderGroupHandleCaptureReplay      Bool32
	rayTracingPipelineShaderGroupHandleCaptureReplayMixed Bool32
	rayTracingPipelineTraceRaysIndirect                   Bool32
	rayTraversalPrimitiveCulling                          Bool32
}

// PhysicalDeviceRayTracingPipelinePropertiesKHR extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceRayTracingPipelinePropertiesKHR = C.VkPhysicalDeviceRayTracingPipelinePropertiesKHR

@[typedef]
pub struct C.VkPhysicalDeviceRayTracingPipelinePropertiesKHR {
pub mut:
	sType                              StructureType = StructureType.physical_device_ray_tracing_pipeline_properties_khr
	pNext                              voidptr       = unsafe { nil }
	shaderGroupHandleSize              u32
	maxRayRecursionDepth               u32
	maxShaderGroupStride               u32
	shaderGroupBaseAlignment           u32
	shaderGroupHandleCaptureReplaySize u32
	maxRayDispatchInvocationCount      u32
	shaderGroupHandleAlignment         u32
	maxRayHitAttributeSize             u32
}

pub type TraceRaysIndirectCommandKHR = C.VkTraceRaysIndirectCommandKHR

@[typedef]
pub struct C.VkTraceRaysIndirectCommandKHR {
pub mut:
	width  u32
	height u32
	depth  u32
}

@[keep_args_alive]
fn C.vkCmdTraceRaysKHR(command_buffer CommandBuffer, p_raygen_shader_binding_table &StridedDeviceAddressRegionKHR, p_miss_shader_binding_table &StridedDeviceAddressRegionKHR, p_hit_shader_binding_table &StridedDeviceAddressRegionKHR, p_callable_shader_binding_table &StridedDeviceAddressRegionKHR, width u32, height u32, depth u32)

pub type PFN_vkCmdTraceRaysKHR = fn (command_buffer CommandBuffer, p_raygen_shader_binding_table &StridedDeviceAddressRegionKHR, p_miss_shader_binding_table &StridedDeviceAddressRegionKHR, p_hit_shader_binding_table &StridedDeviceAddressRegionKHR, p_callable_shader_binding_table &StridedDeviceAddressRegionKHR, width u32, height u32, depth u32)

@[inline]
pub fn cmd_trace_rays_khr(command_buffer CommandBuffer,
	p_raygen_shader_binding_table &StridedDeviceAddressRegionKHR,
	p_miss_shader_binding_table &StridedDeviceAddressRegionKHR,
	p_hit_shader_binding_table &StridedDeviceAddressRegionKHR,
	p_callable_shader_binding_table &StridedDeviceAddressRegionKHR,
	width u32,
	height u32,
	depth u32) {
	C.vkCmdTraceRaysKHR(command_buffer, p_raygen_shader_binding_table, p_miss_shader_binding_table,
		p_hit_shader_binding_table, p_callable_shader_binding_table, width, height, depth)
}

@[keep_args_alive]
fn C.vkCreateRayTracingPipelinesKHR(device Device, deferred_operation DeferredOperationKHR, pipeline_cache PipelineCache, create_info_count u32, p_create_infos &RayTracingPipelineCreateInfoKHR, p_allocator &AllocationCallbacks, p_pipelines &Pipeline) Result

pub type PFN_vkCreateRayTracingPipelinesKHR = fn (device Device, deferred_operation DeferredOperationKHR, pipeline_cache PipelineCache, create_info_count u32, p_create_infos &RayTracingPipelineCreateInfoKHR, p_allocator &AllocationCallbacks, p_pipelines &Pipeline) Result

@[inline]
pub fn create_ray_tracing_pipelines_khr(device Device,
	deferred_operation DeferredOperationKHR,
	pipeline_cache PipelineCache,
	create_info_count u32,
	p_create_infos &RayTracingPipelineCreateInfoKHR,
	p_allocator &AllocationCallbacks,
	p_pipelines &Pipeline) Result {
	return C.vkCreateRayTracingPipelinesKHR(device, deferred_operation, pipeline_cache,
		create_info_count, p_create_infos, p_allocator, p_pipelines)
}

@[keep_args_alive]
fn C.vkGetRayTracingCaptureReplayShaderGroupHandlesKHR(device Device, pipeline Pipeline, first_group u32, group_count u32, data_size usize, p_data voidptr) Result

pub type PFN_vkGetRayTracingCaptureReplayShaderGroupHandlesKHR = fn (device Device, pipeline Pipeline, first_group u32, group_count u32, data_size usize, p_data voidptr) Result

@[inline]
pub fn get_ray_tracing_capture_replay_shader_group_handles_khr(device Device,
	pipeline Pipeline,
	first_group u32,
	group_count u32,
	data_size usize,
	p_data voidptr) Result {
	return C.vkGetRayTracingCaptureReplayShaderGroupHandlesKHR(device, pipeline, first_group,
		group_count, data_size, p_data)
}

@[keep_args_alive]
fn C.vkCmdTraceRaysIndirectKHR(command_buffer CommandBuffer, p_raygen_shader_binding_table &StridedDeviceAddressRegionKHR, p_miss_shader_binding_table &StridedDeviceAddressRegionKHR, p_hit_shader_binding_table &StridedDeviceAddressRegionKHR, p_callable_shader_binding_table &StridedDeviceAddressRegionKHR, indirect_device_address DeviceAddress)

pub type PFN_vkCmdTraceRaysIndirectKHR = fn (command_buffer CommandBuffer, p_raygen_shader_binding_table &StridedDeviceAddressRegionKHR, p_miss_shader_binding_table &StridedDeviceAddressRegionKHR, p_hit_shader_binding_table &StridedDeviceAddressRegionKHR, p_callable_shader_binding_table &StridedDeviceAddressRegionKHR, indirect_device_address DeviceAddress)

@[inline]
pub fn cmd_trace_rays_indirect_khr(command_buffer CommandBuffer,
	p_raygen_shader_binding_table &StridedDeviceAddressRegionKHR,
	p_miss_shader_binding_table &StridedDeviceAddressRegionKHR,
	p_hit_shader_binding_table &StridedDeviceAddressRegionKHR,
	p_callable_shader_binding_table &StridedDeviceAddressRegionKHR,
	indirect_device_address DeviceAddress) {
	C.vkCmdTraceRaysIndirectKHR(command_buffer, p_raygen_shader_binding_table, p_miss_shader_binding_table,
		p_hit_shader_binding_table, p_callable_shader_binding_table, indirect_device_address)
}

@[keep_args_alive]
fn C.vkGetRayTracingShaderGroupStackSizeKHR(device Device, pipeline Pipeline, group u32, group_shader ShaderGroupShaderKHR) DeviceSize

pub type PFN_vkGetRayTracingShaderGroupStackSizeKHR = fn (device Device, pipeline Pipeline, group u32, group_shader ShaderGroupShaderKHR) DeviceSize

@[inline]
pub fn get_ray_tracing_shader_group_stack_size_khr(device Device,
	pipeline Pipeline,
	group u32,
	group_shader ShaderGroupShaderKHR) DeviceSize {
	return C.vkGetRayTracingShaderGroupStackSizeKHR(device, pipeline, group, group_shader)
}

@[keep_args_alive]
fn C.vkCmdSetRayTracingPipelineStackSizeKHR(command_buffer CommandBuffer, pipeline_stack_size u32)

pub type PFN_vkCmdSetRayTracingPipelineStackSizeKHR = fn (command_buffer CommandBuffer, pipeline_stack_size u32)

@[inline]
pub fn cmd_set_ray_tracing_pipeline_stack_size_khr(command_buffer CommandBuffer,
	pipeline_stack_size u32) {
	C.vkCmdSetRayTracingPipelineStackSizeKHR(command_buffer, pipeline_stack_size)
}

pub const khr_ray_query_spec_version = 1
pub const khr_ray_query_extension_name = c'VK_KHR_ray_query'
// PhysicalDeviceRayQueryFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceRayQueryFeaturesKHR = C.VkPhysicalDeviceRayQueryFeaturesKHR

@[typedef]
pub struct C.VkPhysicalDeviceRayQueryFeaturesKHR {
pub mut:
	sType    StructureType = StructureType.physical_device_ray_query_features_khr
	pNext    voidptr       = unsafe { nil }
	rayQuery Bool32
}

pub const ext_mesh_shader_spec_version = 1
pub const ext_mesh_shader_extension_name = c'VK_EXT_mesh_shader'
// PhysicalDeviceMeshShaderFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub type PhysicalDeviceMeshShaderFeaturesEXT = C.VkPhysicalDeviceMeshShaderFeaturesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMeshShaderFeaturesEXT {
pub mut:
	sType                                  StructureType = StructureType.physical_device_mesh_shader_features_ext
	pNext                                  voidptr       = unsafe { nil }
	taskShader                             Bool32
	meshShader                             Bool32
	multiviewMeshShader                    Bool32
	primitiveFragmentShadingRateMeshShader Bool32
	meshShaderQueries                      Bool32
}

// PhysicalDeviceMeshShaderPropertiesEXT extends VkPhysicalDeviceProperties2
pub type PhysicalDeviceMeshShaderPropertiesEXT = C.VkPhysicalDeviceMeshShaderPropertiesEXT

@[typedef]
pub struct C.VkPhysicalDeviceMeshShaderPropertiesEXT {
pub mut:
	sType                                 StructureType = StructureType.physical_device_mesh_shader_properties_ext
	pNext                                 voidptr       = unsafe { nil }
	maxTaskWorkGroupTotalCount            u32
	maxTaskWorkGroupCount                 [3]u32
	maxTaskWorkGroupInvocations           u32
	maxTaskWorkGroupSize                  [3]u32
	maxTaskPayloadSize                    u32
	maxTaskSharedMemorySize               u32
	maxTaskPayloadAndSharedMemorySize     u32
	maxMeshWorkGroupTotalCount            u32
	maxMeshWorkGroupCount                 [3]u32
	maxMeshWorkGroupInvocations           u32
	maxMeshWorkGroupSize                  [3]u32
	maxMeshSharedMemorySize               u32
	maxMeshPayloadAndSharedMemorySize     u32
	maxMeshOutputMemorySize               u32
	maxMeshPayloadAndOutputMemorySize     u32
	maxMeshOutputComponents               u32
	maxMeshOutputVertices                 u32
	maxMeshOutputPrimitives               u32
	maxMeshOutputLayers                   u32
	maxMeshMultiviewViewCount             u32
	meshOutputPerVertexGranularity        u32
	meshOutputPerPrimitiveGranularity     u32
	maxPreferredTaskWorkGroupInvocations  u32
	maxPreferredMeshWorkGroupInvocations  u32
	prefersLocalInvocationVertexOutput    Bool32
	prefersLocalInvocationPrimitiveOutput Bool32
	prefersCompactVertexOutput            Bool32
	prefersCompactPrimitiveOutput         Bool32
}

pub type DrawMeshTasksIndirectCommandEXT = C.VkDrawMeshTasksIndirectCommandEXT

@[typedef]
pub struct C.VkDrawMeshTasksIndirectCommandEXT {
pub mut:
	groupCountX u32
	groupCountY u32
	groupCountZ u32
}

@[keep_args_alive]
fn C.vkCmdDrawMeshTasksEXT(command_buffer CommandBuffer, group_count_x u32, group_count_y u32, group_count_z u32)

pub type PFN_vkCmdDrawMeshTasksEXT = fn (command_buffer CommandBuffer, group_count_x u32, group_count_y u32, group_count_z u32)

@[inline]
pub fn cmd_draw_mesh_tasks_ext(command_buffer CommandBuffer,
	group_count_x u32,
	group_count_y u32,
	group_count_z u32) {
	C.vkCmdDrawMeshTasksEXT(command_buffer, group_count_x, group_count_y, group_count_z)
}

@[keep_args_alive]
fn C.vkCmdDrawMeshTasksIndirectEXT(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, draw_count u32, stride u32)

pub type PFN_vkCmdDrawMeshTasksIndirectEXT = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_mesh_tasks_indirect_ext(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	draw_count u32,
	stride u32) {
	C.vkCmdDrawMeshTasksIndirectEXT(command_buffer, buffer, offset, draw_count, stride)
}

@[keep_args_alive]
fn C.vkCmdDrawMeshTasksIndirectCountEXT(command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

pub type PFN_vkCmdDrawMeshTasksIndirectCountEXT = fn (command_buffer CommandBuffer, buffer Buffer, offset DeviceSize, count_buffer Buffer, count_buffer_offset DeviceSize, max_draw_count u32, stride u32)

@[inline]
pub fn cmd_draw_mesh_tasks_indirect_count_ext(command_buffer CommandBuffer,
	buffer Buffer,
	offset DeviceSize,
	count_buffer Buffer,
	count_buffer_offset DeviceSize,
	max_draw_count u32,
	stride u32) {
	C.vkCmdDrawMeshTasksIndirectCountEXT(command_buffer, buffer, offset, count_buffer,
		count_buffer_offset, max_draw_count, stride)
}
