module vulkan

/*
** Copyright 2024 antono2@github.com.
**
** SPDX-License-Identifier: LGPL-2.1-only
*/

/*
** This module is generated from the Khronos Vulkan XML API Registry.
**
*/

import dl
import dl.loader

#flag -I @VMODROOT/include/vk_video
#include "vulkan_video_codec_h264std.h"
#include "vulkan_video_codec_h264std_decode.h"
#include "vulkan_video_codec_h264std_encode.h"
#include "vulkan_video_codec_h265std.h"
#include "vulkan_video_codec_h265std_decode.h"
#include "vulkan_video_codec_h265std_encode.h"
#include "vulkan_video_codecs_common.h"

@[heap]
const loader_instance = *loader.get_or_create_dynamic_lib_loader(loader.DynamicLibLoaderConfig{
	flags: dl.rtld_lazy
	key: 'vulkan'
	env_path: '' // LD_LIBRARY_PATH environment variable is searched by default
	paths: ['libvulkan.so.1', 'vulkan-1.dll']
}) or { panic("Couldn't create vulkan loader") }
pub const loader_p = &loader_instance


// VK_VERSION_1_0 is a preprocessor guard. Do not pass it to API calls.
const version_1_0 = 1

pub fn make_api_version(variant u32, major u32, minor u32, patch u32) u32 {
  return variant << 29 | major << 22 | minor << 12 | patch
}

pub const api_version_1_0 = make_api_version(0, 1, 0, 0) // Patch version should always be set to 0
pub const header_version = 272

pub const header_version_complete = make_api_version(0, 1, 3, header_version)
pub fn version_variant(version u32) u32 {
  return version >> 29
}
pub fn api_version_major(version u32) u32 {
  return version >> 22 & u32(0x7F)
}
pub fn api_version_minor(version u32) u32 {
  return version >> 12 & u32(0x3FF)
}
pub fn api_version_patch(version u32) u32 {
  return version & u32(0xFFF)
}
pub type Bool32 = u32
pub type DeviceAddress = u64
pub type DeviceSize = u64
pub type Flags = u32
pub type SampleMask = u32
pub type C.Buffer = voidptr
pub type C.Image = voidptr
pub type C.Instance = voidptr
pub type C.PhysicalDevice = voidptr
pub type C.Device = voidptr
pub type C.Queue = voidptr
pub type C.Semaphore = voidptr
pub type C.CommandBuffer = voidptr
pub type C.Fence = voidptr
pub type C.DeviceMemory = voidptr
pub type C.Event = voidptr
pub type C.QueryPool = voidptr
pub type C.BufferView = voidptr
pub type C.ImageView = voidptr
pub type C.ShaderModule = voidptr
pub type C.PipelineCache = voidptr
pub type C.PipelineLayout = voidptr
pub type C.Pipeline = voidptr
pub type C.RenderPass = voidptr
pub type C.DescriptorSetLayout = voidptr
pub type C.Sampler = voidptr
pub type C.DescriptorSet = voidptr
pub type C.DescriptorPool = voidptr
pub type C.Framebuffer = voidptr
pub type C.CommandPool = voidptr
pub const attachment_unused                 = ~u32(0)
pub const vk_false                          = u32(0)
pub const lod_clamp_none                    = f32(1000.0)
pub const queue_family_ignored              = ~u32(0)
pub const remaining_array_layers            = ~u32(0)
pub const remaining_mip_levels              = ~u32(0)
pub const subpass_external                  = ~u32(0)
pub const vk_true                           = u32(1)
pub const whole_size                        = ~u64(0)
pub const max_memory_types                  = u32(32)
pub const max_physical_device_name_size     = u32(256)
pub const uuid_size                         = u32(16)
pub const max_extension_name_size           = u32(256)
pub const max_description_size              = u32(256)
pub const max_memory_heaps                  = u32(16)

pub enum Result {
    success = int(0)
    not_ready = int(1)
    timeout = int(2)
    event_set = int(3)
    event_reset = int(4)
    incomplete = int(5)
    error_out_of_host_memory = int(-1)
    error_out_of_device_memory = int(-2)
    error_initialization_failed = int(-3)
    error_device_lost = int(-4)
    error_memory_map_failed = int(-5)
    error_layer_not_present = int(-6)
    error_extension_not_present = int(-7)
    error_feature_not_present = int(-8)
    error_incompatible_driver = int(-9)
    error_too_many_objects = int(-10)
    error_format_not_supported = int(-11)
    error_fragmented_pool = int(-12)
    error_unknown = int(-13)
    error_out_of_pool_memory = int(-1000069000)
    error_invalid_external_handle = int(-1000072003)
    error_fragmentation = int(-1000161000)
    error_invalid_opaque_capture_address = int(-1000257000)
    pipeline_compile_required = int(1000297000)
    error_surface_lost_khr = int(-1000000000)
    error_native_window_in_use_khr = int(-1000000001)
    suboptimal_khr = int(1000001003)
    error_out_of_date_khr = int(-1000001004)
    error_incompatible_display_khr = int(-1000003001)
    error_validation_failed_ext = int(-1000011001)
    error_invalid_shader_nv = int(-1000012000)
    error_image_usage_not_supported_khr = int(-1000023000)
    error_video_picture_layout_not_supported_khr = int(-1000023001)
    error_video_profile_operation_not_supported_khr = int(-1000023002)
    error_video_profile_format_not_supported_khr = int(-1000023003)
    error_video_profile_codec_not_supported_khr = int(-1000023004)
    error_video_std_version_not_supported_khr = int(-1000023005)
    error_invalid_drm_format_modifier_plane_layout_ext = int(-1000158000)
    error_not_permitted_khr = int(-1000174001)
    error_full_screen_exclusive_mode_lost_ext = int(-1000255000)
    thread_idle_khr = int(1000268000)
    thread_done_khr = int(1000268001)
    operation_deferred_khr = int(1000268002)
    operation_not_deferred_khr = int(1000268003)
    error_compression_exhausted_ext = int(-1000338000)
    error_incompatible_shader_binary_ext = int(1000482000)
    result_max_enum = int(0x7FFFFFFF)
}


pub enum StructureType {
    structure_type_application_info = int(0)
    structure_type_instance_create_info = int(1)
    structure_type_device_queue_create_info = int(2)
    structure_type_device_create_info = int(3)
    structure_type_submit_info = int(4)
    structure_type_memory_allocate_info = int(5)
    structure_type_mapped_memory_range = int(6)
    structure_type_bind_sparse_info = int(7)
    structure_type_fence_create_info = int(8)
    structure_type_semaphore_create_info = int(9)
    structure_type_event_create_info = int(10)
    structure_type_query_pool_create_info = int(11)
    structure_type_buffer_create_info = int(12)
    structure_type_buffer_view_create_info = int(13)
    structure_type_image_create_info = int(14)
    structure_type_image_view_create_info = int(15)
    structure_type_shader_module_create_info = int(16)
    structure_type_pipeline_cache_create_info = int(17)
    structure_type_pipeline_shader_stage_create_info = int(18)
    structure_type_pipeline_vertex_input_state_create_info = int(19)
    structure_type_pipeline_input_assembly_state_create_info = int(20)
    structure_type_pipeline_tessellation_state_create_info = int(21)
    structure_type_pipeline_viewport_state_create_info = int(22)
    structure_type_pipeline_rasterization_state_create_info = int(23)
    structure_type_pipeline_multisample_state_create_info = int(24)
    structure_type_pipeline_depth_stencil_state_create_info = int(25)
    structure_type_pipeline_color_blend_state_create_info = int(26)
    structure_type_pipeline_dynamic_state_create_info = int(27)
    structure_type_graphics_pipeline_create_info = int(28)
    structure_type_compute_pipeline_create_info = int(29)
    structure_type_pipeline_layout_create_info = int(30)
    structure_type_sampler_create_info = int(31)
    structure_type_descriptor_set_layout_create_info = int(32)
    structure_type_descriptor_pool_create_info = int(33)
    structure_type_descriptor_set_allocate_info = int(34)
    structure_type_write_descriptor_set = int(35)
    structure_type_copy_descriptor_set = int(36)
    structure_type_framebuffer_create_info = int(37)
    structure_type_render_pass_create_info = int(38)
    structure_type_command_pool_create_info = int(39)
    structure_type_command_buffer_allocate_info = int(40)
    structure_type_command_buffer_inheritance_info = int(41)
    structure_type_command_buffer_begin_info = int(42)
    structure_type_render_pass_begin_info = int(43)
    structure_type_buffer_memory_barrier = int(44)
    structure_type_image_memory_barrier = int(45)
    structure_type_memory_barrier = int(46)
    structure_type_loader_instance_create_info = int(47)
    structure_type_loader_device_create_info = int(48)
    structure_type_physical_device_subgroup_properties = int(1000094000)
    structure_type_bind_buffer_memory_info = int(1000157000)
    structure_type_bind_image_memory_info = int(1000157001)
    structure_type_physical_device_16bit_storage_features = int(1000083000)
    structure_type_memory_dedicated_requirements = int(1000127000)
    structure_type_memory_dedicated_allocate_info = int(1000127001)
    structure_type_memory_allocate_flags_info = int(1000060000)
    structure_type_device_group_render_pass_begin_info = int(1000060003)
    structure_type_device_group_command_buffer_begin_info = int(1000060004)
    structure_type_device_group_submit_info = int(1000060005)
    structure_type_device_group_bind_sparse_info = int(1000060006)
    structure_type_bind_buffer_memory_device_group_info = int(1000060013)
    structure_type_bind_image_memory_device_group_info = int(1000060014)
    structure_type_physical_device_group_properties = int(1000070000)
    structure_type_device_group_device_create_info = int(1000070001)
    structure_type_buffer_memory_requirements_info_2 = int(1000146000)
    structure_type_image_memory_requirements_info_2 = int(1000146001)
    structure_type_image_sparse_memory_requirements_info_2 = int(1000146002)
    structure_type_memory_requirements_2 = int(1000146003)
    structure_type_sparse_image_memory_requirements_2 = int(1000146004)
    structure_type_physical_device_features_2 = int(1000059000)
    structure_type_physical_device_properties_2 = int(1000059001)
    structure_type_format_properties_2 = int(1000059002)
    structure_type_image_format_properties_2 = int(1000059003)
    structure_type_physical_device_image_format_info_2 = int(1000059004)
    structure_type_queue_family_properties_2 = int(1000059005)
    structure_type_physical_device_memory_properties_2 = int(1000059006)
    structure_type_sparse_image_format_properties_2 = int(1000059007)
    structure_type_physical_device_sparse_image_format_info_2 = int(1000059008)
    structure_type_physical_device_point_clipping_properties = int(1000117000)
    structure_type_render_pass_input_attachment_aspect_create_info = int(1000117001)
    structure_type_image_view_usage_create_info = int(1000117002)
    structure_type_pipeline_tessellation_domain_origin_state_create_info = int(1000117003)
    structure_type_render_pass_multiview_create_info = int(1000053000)
    structure_type_physical_device_multiview_features = int(1000053001)
    structure_type_physical_device_multiview_properties = int(1000053002)
    structure_type_physical_device_variable_pointers_features = int(1000120000)
    structure_type_protected_submit_info = int(1000145000)
    structure_type_physical_device_protected_memory_features = int(1000145001)
    structure_type_physical_device_protected_memory_properties = int(1000145002)
    structure_type_device_queue_info_2 = int(1000145003)
    structure_type_sampler_ycbcr_conversion_create_info = int(1000156000)
    structure_type_sampler_ycbcr_conversion_info = int(1000156001)
    structure_type_bind_image_plane_memory_info = int(1000156002)
    structure_type_image_plane_memory_requirements_info = int(1000156003)
    structure_type_physical_device_sampler_ycbcr_conversion_features = int(1000156004)
    structure_type_sampler_ycbcr_conversion_image_format_properties = int(1000156005)
    structure_type_descriptor_update_template_create_info = int(1000085000)
    structure_type_physical_device_external_image_format_info = int(1000071000)
    structure_type_external_image_format_properties = int(1000071001)
    structure_type_physical_device_external_buffer_info = int(1000071002)
    structure_type_external_buffer_properties = int(1000071003)
    structure_type_physical_device_id_properties = int(1000071004)
    structure_type_external_memory_buffer_create_info = int(1000072000)
    structure_type_external_memory_image_create_info = int(1000072001)
    structure_type_export_memory_allocate_info = int(1000072002)
    structure_type_physical_device_external_fence_info = int(1000112000)
    structure_type_external_fence_properties = int(1000112001)
    structure_type_export_fence_create_info = int(1000113000)
    structure_type_export_semaphore_create_info = int(1000077000)
    structure_type_physical_device_external_semaphore_info = int(1000076000)
    structure_type_external_semaphore_properties = int(1000076001)
    structure_type_physical_device_maintenance_3_properties = int(1000168000)
    structure_type_descriptor_set_layout_support = int(1000168001)
    structure_type_physical_device_shader_draw_parameters_features = int(1000063000)
    structure_type_physical_device_vulkan_1_1_features = int(49)
    structure_type_physical_device_vulkan_1_1_properties = int(50)
    structure_type_physical_device_vulkan_1_2_features = int(51)
    structure_type_physical_device_vulkan_1_2_properties = int(52)
    structure_type_image_format_list_create_info = int(1000147000)
    structure_type_attachment_description_2 = int(1000109000)
    structure_type_attachment_reference_2 = int(1000109001)
    structure_type_subpass_description_2 = int(1000109002)
    structure_type_subpass_dependency_2 = int(1000109003)
    structure_type_render_pass_create_info_2 = int(1000109004)
    structure_type_subpass_begin_info = int(1000109005)
    structure_type_subpass_end_info = int(1000109006)
    structure_type_physical_device_8bit_storage_features = int(1000177000)
    structure_type_physical_device_driver_properties = int(1000196000)
    structure_type_physical_device_shader_atomic_int64_features = int(1000180000)
    structure_type_physical_device_shader_float16_int8_features = int(1000082000)
    structure_type_physical_device_float_controls_properties = int(1000197000)
    structure_type_descriptor_set_layout_binding_flags_create_info = int(1000161000)
    structure_type_physical_device_descriptor_indexing_features = int(1000161001)
    structure_type_physical_device_descriptor_indexing_properties = int(1000161002)
    structure_type_descriptor_set_variable_descriptor_count_allocate_info = int(1000161003)
    structure_type_descriptor_set_variable_descriptor_count_layout_support = int(1000161004)
    structure_type_physical_device_depth_stencil_resolve_properties = int(1000199000)
    structure_type_subpass_description_depth_stencil_resolve = int(1000199001)
    structure_type_physical_device_scalar_block_layout_features = int(1000221000)
    structure_type_image_stencil_usage_create_info = int(1000246000)
    structure_type_physical_device_sampler_filter_minmax_properties = int(1000130000)
    structure_type_sampler_reduction_mode_create_info = int(1000130001)
    structure_type_physical_device_vulkan_memory_model_features = int(1000211000)
    structure_type_physical_device_imageless_framebuffer_features = int(1000108000)
    structure_type_framebuffer_attachments_create_info = int(1000108001)
    structure_type_framebuffer_attachment_image_info = int(1000108002)
    structure_type_render_pass_attachment_begin_info = int(1000108003)
    structure_type_physical_device_uniform_buffer_standard_layout_features = int(1000253000)
    structure_type_physical_device_shader_subgroup_extended_types_features = int(1000175000)
    structure_type_physical_device_separate_depth_stencil_layouts_features = int(1000241000)
    structure_type_attachment_reference_stencil_layout = int(1000241001)
    structure_type_attachment_description_stencil_layout = int(1000241002)
    structure_type_physical_device_host_query_reset_features = int(1000261000)
    structure_type_physical_device_timeline_semaphore_features = int(1000207000)
    structure_type_physical_device_timeline_semaphore_properties = int(1000207001)
    structure_type_semaphore_type_create_info = int(1000207002)
    structure_type_timeline_semaphore_submit_info = int(1000207003)
    structure_type_semaphore_wait_info = int(1000207004)
    structure_type_semaphore_signal_info = int(1000207005)
    structure_type_physical_device_buffer_device_address_features = int(1000257000)
    structure_type_buffer_device_address_info = int(1000244001)
    structure_type_buffer_opaque_capture_address_create_info = int(1000257002)
    structure_type_memory_opaque_capture_address_allocate_info = int(1000257003)
    structure_type_device_memory_opaque_capture_address_info = int(1000257004)
    structure_type_physical_device_vulkan_1_3_features = int(53)
    structure_type_physical_device_vulkan_1_3_properties = int(54)
    structure_type_pipeline_creation_feedback_create_info = int(1000192000)
    structure_type_physical_device_shader_terminate_invocation_features = int(1000215000)
    structure_type_physical_device_tool_properties = int(1000245000)
    structure_type_physical_device_shader_demote_to_helper_invocation_features = int(1000276000)
    structure_type_physical_device_private_data_features = int(1000295000)
    structure_type_device_private_data_create_info = int(1000295001)
    structure_type_private_data_slot_create_info = int(1000295002)
    structure_type_physical_device_pipeline_creation_cache_control_features = int(1000297000)
    structure_type_memory_barrier_2 = int(1000314000)
    structure_type_buffer_memory_barrier_2 = int(1000314001)
    structure_type_image_memory_barrier_2 = int(1000314002)
    structure_type_dependency_info = int(1000314003)
    structure_type_submit_info_2 = int(1000314004)
    structure_type_semaphore_submit_info = int(1000314005)
    structure_type_command_buffer_submit_info = int(1000314006)
    structure_type_physical_device_synchronization_2_features = int(1000314007)
    structure_type_physical_device_zero_initialize_workgroup_memory_features = int(1000325000)
    structure_type_physical_device_image_robustness_features = int(1000335000)
    structure_type_copy_buffer_info_2 = int(1000337000)
    structure_type_copy_image_info_2 = int(1000337001)
    structure_type_copy_buffer_to_image_info_2 = int(1000337002)
    structure_type_copy_image_to_buffer_info_2 = int(1000337003)
    structure_type_blit_image_info_2 = int(1000337004)
    structure_type_resolve_image_info_2 = int(1000337005)
    structure_type_buffer_copy_2 = int(1000337006)
    structure_type_image_copy_2 = int(1000337007)
    structure_type_image_blit_2 = int(1000337008)
    structure_type_buffer_image_copy_2 = int(1000337009)
    structure_type_image_resolve_2 = int(1000337010)
    structure_type_physical_device_subgroup_size_control_properties = int(1000225000)
    structure_type_pipeline_shader_stage_required_subgroup_size_create_info = int(1000225001)
    structure_type_physical_device_subgroup_size_control_features = int(1000225002)
    structure_type_physical_device_inline_uniform_block_features = int(1000138000)
    structure_type_physical_device_inline_uniform_block_properties = int(1000138001)
    structure_type_write_descriptor_set_inline_uniform_block = int(1000138002)
    structure_type_descriptor_pool_inline_uniform_block_create_info = int(1000138003)
    structure_type_physical_device_texture_compression_astc_hdr_features = int(1000066000)
    structure_type_rendering_info = int(1000044000)
    structure_type_rendering_attachment_info = int(1000044001)
    structure_type_pipeline_rendering_create_info = int(1000044002)
    structure_type_physical_device_dynamic_rendering_features = int(1000044003)
    structure_type_command_buffer_inheritance_rendering_info = int(1000044004)
    structure_type_physical_device_shader_integer_dot_product_features = int(1000280000)
    structure_type_physical_device_shader_integer_dot_product_properties = int(1000280001)
    structure_type_physical_device_texel_buffer_alignment_properties = int(1000281001)
    structure_type_format_properties_3 = int(1000360000)
    structure_type_physical_device_maintenance_4_features = int(1000413000)
    structure_type_physical_device_maintenance_4_properties = int(1000413001)
    structure_type_device_buffer_memory_requirements = int(1000413002)
    structure_type_device_image_memory_requirements = int(1000413003)
    structure_type_swapchain_create_info_khr = int(1000001000)
    structure_type_present_info_khr = int(1000001001)
    structure_type_device_group_present_capabilities_khr = int(1000060007)
    structure_type_image_swapchain_create_info_khr = int(1000060008)
    structure_type_bind_image_memory_swapchain_info_khr = int(1000060009)
    structure_type_acquire_next_image_info_khr = int(1000060010)
    structure_type_device_group_present_info_khr = int(1000060011)
    structure_type_device_group_swapchain_create_info_khr = int(1000060012)
    structure_type_display_mode_create_info_khr = int(1000002000)
    structure_type_display_surface_create_info_khr = int(1000002001)
    structure_type_display_present_info_khr = int(1000003000)
    structure_type_xlib_surface_create_info_khr = int(1000004000)
    structure_type_xcb_surface_create_info_khr = int(1000005000)
    structure_type_wayland_surface_create_info_khr = int(1000006000)
    structure_type_android_surface_create_info_khr = int(1000008000)
    structure_type_win32_surface_create_info_khr = int(1000009000)
    structure_type_debug_report_callback_create_info_ext = int(1000011000)
    structure_type_pipeline_rasterization_state_rasterization_order_amd = int(1000018000)
    structure_type_debug_marker_object_name_info_ext = int(1000022000)
    structure_type_debug_marker_object_tag_info_ext = int(1000022001)
    structure_type_debug_marker_marker_info_ext = int(1000022002)
    structure_type_video_profile_info_khr = int(1000023000)
    structure_type_video_capabilities_khr = int(1000023001)
    structure_type_video_picture_resource_info_khr = int(1000023002)
    structure_type_video_session_memory_requirements_khr = int(1000023003)
    structure_type_bind_video_session_memory_info_khr = int(1000023004)
    structure_type_video_session_create_info_khr = int(1000023005)
    structure_type_video_session_parameters_create_info_khr = int(1000023006)
    structure_type_video_session_parameters_update_info_khr = int(1000023007)
    structure_type_video_begin_coding_info_khr = int(1000023008)
    structure_type_video_end_coding_info_khr = int(1000023009)
    structure_type_video_coding_control_info_khr = int(1000023010)
    structure_type_video_reference_slot_info_khr = int(1000023011)
    structure_type_queue_family_video_properties_khr = int(1000023012)
    structure_type_video_profile_list_info_khr = int(1000023013)
    structure_type_physical_device_video_format_info_khr = int(1000023014)
    structure_type_video_format_properties_khr = int(1000023015)
    structure_type_queue_family_query_result_status_properties_khr = int(1000023016)
    structure_type_video_decode_info_khr = int(1000024000)
    structure_type_video_decode_capabilities_khr = int(1000024001)
    structure_type_video_decode_usage_info_khr = int(1000024002)
    structure_type_dedicated_allocation_image_create_info_nv = int(1000026000)
    structure_type_dedicated_allocation_buffer_create_info_nv = int(1000026001)
    structure_type_dedicated_allocation_memory_allocate_info_nv = int(1000026002)
    structure_type_physical_device_transform_feedback_features_ext = int(1000028000)
    structure_type_physical_device_transform_feedback_properties_ext = int(1000028001)
    structure_type_pipeline_rasterization_state_stream_create_info_ext = int(1000028002)
    structure_type_cu_module_create_info_nvx = int(1000029000)
    structure_type_cu_function_create_info_nvx = int(1000029001)
    structure_type_cu_launch_info_nvx = int(1000029002)
    structure_type_image_view_handle_info_nvx = int(1000030000)
    structure_type_image_view_address_properties_nvx = int(1000030001)
    structure_type_video_decode_h264_capabilities_khr = int(1000040000)
    structure_type_video_decode_h264_picture_info_khr = int(1000040001)
    structure_type_video_decode_h264_profile_info_khr = int(1000040003)
    structure_type_video_decode_h264_session_parameters_create_info_khr = int(1000040004)
    structure_type_video_decode_h264_session_parameters_add_info_khr = int(1000040005)
    structure_type_video_decode_h264_dpb_slot_info_khr = int(1000040006)
    structure_type_texture_lod_gather_format_properties_amd = int(1000041000)
    structure_type_rendering_fragment_shading_rate_attachment_info_khr = int(1000044006)
    structure_type_rendering_fragment_density_map_attachment_info_ext = int(1000044007)
    structure_type_attachment_sample_count_info_amd = int(1000044008)
    structure_type_multiview_per_view_attributes_info_nvx = int(1000044009)
    structure_type_stream_descriptor_surface_create_info_ggp = int(1000049000)
    structure_type_physical_device_corner_sampled_image_features_nv = int(1000050000)
    structure_type_external_memory_image_create_info_nv = int(1000056000)
    structure_type_export_memory_allocate_info_nv = int(1000056001)
    structure_type_import_memory_win32_handle_info_nv = int(1000057000)
    structure_type_export_memory_win32_handle_info_nv = int(1000057001)
    structure_type_win32_keyed_mutex_acquire_release_info_nv = int(1000058000)
    structure_type_validation_flags_ext = int(1000061000)
    structure_type_vi_surface_create_info_nn = int(1000062000)
    structure_type_image_view_astc_decode_mode_ext = int(1000067000)
    structure_type_physical_device_astc_decode_features_ext = int(1000067001)
    structure_type_pipeline_robustness_create_info_ext = int(1000068000)
    structure_type_physical_device_pipeline_robustness_features_ext = int(1000068001)
    structure_type_physical_device_pipeline_robustness_properties_ext = int(1000068002)
    structure_type_import_memory_win32_handle_info_khr = int(1000073000)
    structure_type_export_memory_win32_handle_info_khr = int(1000073001)
    structure_type_memory_win32_handle_properties_khr = int(1000073002)
    structure_type_memory_get_win32_handle_info_khr = int(1000073003)
    structure_type_import_memory_fd_info_khr = int(1000074000)
    structure_type_memory_fd_properties_khr = int(1000074001)
    structure_type_memory_get_fd_info_khr = int(1000074002)
    structure_type_win32_keyed_mutex_acquire_release_info_khr = int(1000075000)
    structure_type_import_semaphore_win32_handle_info_khr = int(1000078000)
    structure_type_export_semaphore_win32_handle_info_khr = int(1000078001)
    structure_type_d3d12_fence_submit_info_khr = int(1000078002)
    structure_type_semaphore_get_win32_handle_info_khr = int(1000078003)
    structure_type_import_semaphore_fd_info_khr = int(1000079000)
    structure_type_semaphore_get_fd_info_khr = int(1000079001)
    structure_type_physical_device_push_descriptor_properties_khr = int(1000080000)
    structure_type_command_buffer_inheritance_conditional_rendering_info_ext = int(1000081000)
    structure_type_physical_device_conditional_rendering_features_ext = int(1000081001)
    structure_type_conditional_rendering_begin_info_ext = int(1000081002)
    structure_type_present_regions_khr = int(1000084000)
    structure_type_pipeline_viewport_w_scaling_state_create_info_nv = int(1000087000)
    structure_type_surface_capabilities_2_ext = int(1000090000)
    structure_type_display_power_info_ext = int(1000091000)
    structure_type_device_event_info_ext = int(1000091001)
    structure_type_display_event_info_ext = int(1000091002)
    structure_type_swapchain_counter_create_info_ext = int(1000091003)
    structure_type_present_times_info_google = int(1000092000)
    structure_type_physical_device_multiview_per_view_attributes_properties_nvx = int(1000097000)
    structure_type_pipeline_viewport_swizzle_state_create_info_nv = int(1000098000)
    structure_type_physical_device_discard_rectangle_properties_ext = int(1000099000)
    structure_type_pipeline_discard_rectangle_state_create_info_ext = int(1000099001)
    structure_type_physical_device_conservative_rasterization_properties_ext = int(1000101000)
    structure_type_pipeline_rasterization_conservative_state_create_info_ext = int(1000101001)
    structure_type_physical_device_depth_clip_enable_features_ext = int(1000102000)
    structure_type_pipeline_rasterization_depth_clip_state_create_info_ext = int(1000102001)
    structure_type_hdr_metadata_ext = int(1000105000)
    structure_type_physical_device_relaxed_line_rasterization_features_img = int(1000110000)
    structure_type_shared_present_surface_capabilities_khr = int(1000111000)
    structure_type_import_fence_win32_handle_info_khr = int(1000114000)
    structure_type_export_fence_win32_handle_info_khr = int(1000114001)
    structure_type_fence_get_win32_handle_info_khr = int(1000114002)
    structure_type_import_fence_fd_info_khr = int(1000115000)
    structure_type_fence_get_fd_info_khr = int(1000115001)
    structure_type_physical_device_performance_query_features_khr = int(1000116000)
    structure_type_physical_device_performance_query_properties_khr = int(1000116001)
    structure_type_query_pool_performance_create_info_khr = int(1000116002)
    structure_type_performance_query_submit_info_khr = int(1000116003)
    structure_type_acquire_profiling_lock_info_khr = int(1000116004)
    structure_type_performance_counter_khr = int(1000116005)
    structure_type_performance_counter_description_khr = int(1000116006)
    structure_type_physical_device_surface_info_2_khr = int(1000119000)
    structure_type_surface_capabilities_2_khr = int(1000119001)
    structure_type_surface_format_2_khr = int(1000119002)
    structure_type_display_properties_2_khr = int(1000121000)
    structure_type_display_plane_properties_2_khr = int(1000121001)
    structure_type_display_mode_properties_2_khr = int(1000121002)
    structure_type_display_plane_info_2_khr = int(1000121003)
    structure_type_display_plane_capabilities_2_khr = int(1000121004)
    structure_type_ios_surface_create_info_mvk = int(1000122000)
    structure_type_macos_surface_create_info_mvk = int(1000123000)
    structure_type_debug_utils_object_name_info_ext = int(1000128000)
    structure_type_debug_utils_object_tag_info_ext = int(1000128001)
    structure_type_debug_utils_label_ext = int(1000128002)
    structure_type_debug_utils_messenger_callback_data_ext = int(1000128003)
    structure_type_debug_utils_messenger_create_info_ext = int(1000128004)
    structure_type_android_hardware_buffer_usage_android = int(1000129000)
    structure_type_android_hardware_buffer_properties_android = int(1000129001)
    structure_type_android_hardware_buffer_format_properties_android = int(1000129002)
    structure_type_import_android_hardware_buffer_info_android = int(1000129003)
    structure_type_memory_get_android_hardware_buffer_info_android = int(1000129004)
    structure_type_external_format_android = int(1000129005)
    structure_type_android_hardware_buffer_format_properties_2_android = int(1000129006)
    structure_type_sample_locations_info_ext = int(1000143000)
    structure_type_render_pass_sample_locations_begin_info_ext = int(1000143001)
    structure_type_pipeline_sample_locations_state_create_info_ext = int(1000143002)
    structure_type_physical_device_sample_locations_properties_ext = int(1000143003)
    structure_type_multisample_properties_ext = int(1000143004)
    structure_type_physical_device_blend_operation_advanced_features_ext = int(1000148000)
    structure_type_physical_device_blend_operation_advanced_properties_ext = int(1000148001)
    structure_type_pipeline_color_blend_advanced_state_create_info_ext = int(1000148002)
    structure_type_pipeline_coverage_to_color_state_create_info_nv = int(1000149000)
    structure_type_write_descriptor_set_acceleration_structure_khr = int(1000150007)
    structure_type_acceleration_structure_build_geometry_info_khr = int(1000150000)
    structure_type_acceleration_structure_device_address_info_khr = int(1000150002)
    structure_type_acceleration_structure_geometry_aabbs_data_khr = int(1000150003)
    structure_type_acceleration_structure_geometry_instances_data_khr = int(1000150004)
    structure_type_acceleration_structure_geometry_triangles_data_khr = int(1000150005)
    structure_type_acceleration_structure_geometry_khr = int(1000150006)
    structure_type_acceleration_structure_version_info_khr = int(1000150009)
    structure_type_copy_acceleration_structure_info_khr = int(1000150010)
    structure_type_copy_acceleration_structure_to_memory_info_khr = int(1000150011)
    structure_type_copy_memory_to_acceleration_structure_info_khr = int(1000150012)
    structure_type_physical_device_acceleration_structure_features_khr = int(1000150013)
    structure_type_physical_device_acceleration_structure_properties_khr = int(1000150014)
    structure_type_acceleration_structure_create_info_khr = int(1000150017)
    structure_type_acceleration_structure_build_sizes_info_khr = int(1000150020)
    structure_type_physical_device_ray_tracing_pipeline_features_khr = int(1000347000)
    structure_type_physical_device_ray_tracing_pipeline_properties_khr = int(1000347001)
    structure_type_ray_tracing_pipeline_create_info_khr = int(1000150015)
    structure_type_ray_tracing_shader_group_create_info_khr = int(1000150016)
    structure_type_ray_tracing_pipeline_interface_create_info_khr = int(1000150018)
    structure_type_physical_device_ray_query_features_khr = int(1000348013)
    structure_type_pipeline_coverage_modulation_state_create_info_nv = int(1000152000)
    structure_type_physical_device_shader_sm_builtins_features_nv = int(1000154000)
    structure_type_physical_device_shader_sm_builtins_properties_nv = int(1000154001)
    structure_type_drm_format_modifier_properties_list_ext = int(1000158000)
    structure_type_physical_device_image_drm_format_modifier_info_ext = int(1000158002)
    structure_type_image_drm_format_modifier_list_create_info_ext = int(1000158003)
    structure_type_image_drm_format_modifier_explicit_create_info_ext = int(1000158004)
    structure_type_image_drm_format_modifier_properties_ext = int(1000158005)
    structure_type_drm_format_modifier_properties_list_2_ext = int(1000158006)
    structure_type_validation_cache_create_info_ext = int(1000160000)
    structure_type_shader_module_validation_cache_create_info_ext = int(1000160001)
    structure_type_pipeline_viewport_shading_rate_image_state_create_info_nv = int(1000164000)
    structure_type_physical_device_shading_rate_image_features_nv = int(1000164001)
    structure_type_physical_device_shading_rate_image_properties_nv = int(1000164002)
    structure_type_pipeline_viewport_coarse_sample_order_state_create_info_nv = int(1000164005)
    structure_type_ray_tracing_pipeline_create_info_nv = int(1000165000)
    structure_type_acceleration_structure_create_info_nv = int(1000165001)
    structure_type_geometry_nv = int(1000165003)
    structure_type_geometry_triangles_nv = int(1000165004)
    structure_type_geometry_aabb_nv = int(1000165005)
    structure_type_bind_acceleration_structure_memory_info_nv = int(1000165006)
    structure_type_write_descriptor_set_acceleration_structure_nv = int(1000165007)
    structure_type_acceleration_structure_memory_requirements_info_nv = int(1000165008)
    structure_type_physical_device_ray_tracing_properties_nv = int(1000165009)
    structure_type_ray_tracing_shader_group_create_info_nv = int(1000165011)
    structure_type_acceleration_structure_info_nv = int(1000165012)
    structure_type_physical_device_representative_fragment_test_features_nv = int(1000166000)
    structure_type_pipeline_representative_fragment_test_state_create_info_nv = int(1000166001)
    structure_type_physical_device_image_view_image_format_info_ext = int(1000170000)
    structure_type_filter_cubic_image_view_image_format_properties_ext = int(1000170001)
    structure_type_import_memory_host_pointer_info_ext = int(1000178000)
    structure_type_memory_host_pointer_properties_ext = int(1000178001)
    structure_type_physical_device_external_memory_host_properties_ext = int(1000178002)
    structure_type_physical_device_shader_clock_features_khr = int(1000181000)
    structure_type_pipeline_compiler_control_create_info_amd = int(1000183000)
    structure_type_calibrated_timestamp_info_ext = int(1000184000)
    structure_type_physical_device_shader_core_properties_amd = int(1000185000)
    structure_type_video_decode_h265_capabilities_khr = int(1000187000)
    structure_type_video_decode_h265_session_parameters_create_info_khr = int(1000187001)
    structure_type_video_decode_h265_session_parameters_add_info_khr = int(1000187002)
    structure_type_video_decode_h265_profile_info_khr = int(1000187003)
    structure_type_video_decode_h265_picture_info_khr = int(1000187004)
    structure_type_video_decode_h265_dpb_slot_info_khr = int(1000187005)
    structure_type_device_queue_global_priority_create_info_khr = int(1000174000)
    structure_type_physical_device_global_priority_query_features_khr = int(1000388000)
    structure_type_queue_family_global_priority_properties_khr = int(1000388001)
    structure_type_device_memory_overallocation_create_info_amd = int(1000189000)
    structure_type_physical_device_vertex_attribute_divisor_properties_ext = int(1000190000)
    structure_type_pipeline_vertex_input_divisor_state_create_info_ext = int(1000190001)
    structure_type_physical_device_vertex_attribute_divisor_features_ext = int(1000190002)
    structure_type_present_frame_token_ggp = int(1000191000)
    structure_type_physical_device_compute_shader_derivatives_features_nv = int(1000201000)
    structure_type_physical_device_mesh_shader_features_nv = int(1000202000)
    structure_type_physical_device_mesh_shader_properties_nv = int(1000202001)
    structure_type_physical_device_shader_image_footprint_features_nv = int(1000204000)
    structure_type_pipeline_viewport_exclusive_scissor_state_create_info_nv = int(1000205000)
    structure_type_physical_device_exclusive_scissor_features_nv = int(1000205002)
    structure_type_checkpoint_data_nv = int(1000206000)
    structure_type_queue_family_checkpoint_properties_nv = int(1000206001)
    structure_type_physical_device_shader_integer_functions_2_features_intel = int(1000209000)
    structure_type_query_pool_performance_query_create_info_intel = int(1000210000)
    structure_type_initialize_performance_api_info_intel = int(1000210001)
    structure_type_performance_marker_info_intel = int(1000210002)
    structure_type_performance_stream_marker_info_intel = int(1000210003)
    structure_type_performance_override_info_intel = int(1000210004)
    structure_type_performance_configuration_acquire_info_intel = int(1000210005)
    structure_type_physical_device_pci_bus_info_properties_ext = int(1000212000)
    structure_type_display_native_hdr_surface_capabilities_amd = int(1000213000)
    structure_type_swapchain_display_native_hdr_create_info_amd = int(1000213001)
    structure_type_imagepipe_surface_create_info_fuchsia = int(1000214000)
    structure_type_metal_surface_create_info_ext = int(1000217000)
    structure_type_physical_device_fragment_density_map_features_ext = int(1000218000)
    structure_type_physical_device_fragment_density_map_properties_ext = int(1000218001)
    structure_type_render_pass_fragment_density_map_create_info_ext = int(1000218002)
    structure_type_fragment_shading_rate_attachment_info_khr = int(1000226000)
    structure_type_pipeline_fragment_shading_rate_state_create_info_khr = int(1000226001)
    structure_type_physical_device_fragment_shading_rate_properties_khr = int(1000226002)
    structure_type_physical_device_fragment_shading_rate_features_khr = int(1000226003)
    structure_type_physical_device_fragment_shading_rate_khr = int(1000226004)
    structure_type_physical_device_shader_core_properties_2_amd = int(1000227000)
    structure_type_physical_device_coherent_memory_features_amd = int(1000229000)
    structure_type_physical_device_shader_image_atomic_int64_features_ext = int(1000234000)
    structure_type_physical_device_memory_budget_properties_ext = int(1000237000)
    structure_type_physical_device_memory_priority_features_ext = int(1000238000)
    structure_type_memory_priority_allocate_info_ext = int(1000238001)
    structure_type_surface_protected_capabilities_khr = int(1000239000)
    structure_type_physical_device_dedicated_allocation_image_aliasing_features_nv = int(1000240000)
    structure_type_physical_device_buffer_device_address_features_ext = int(1000244000)
    structure_type_buffer_device_address_create_info_ext = int(1000244002)
    structure_type_validation_features_ext = int(1000247000)
    structure_type_physical_device_present_wait_features_khr = int(1000248000)
    structure_type_physical_device_cooperative_matrix_features_nv = int(1000249000)
    structure_type_cooperative_matrix_properties_nv = int(1000249001)
    structure_type_physical_device_cooperative_matrix_properties_nv = int(1000249002)
    structure_type_physical_device_coverage_reduction_mode_features_nv = int(1000250000)
    structure_type_pipeline_coverage_reduction_state_create_info_nv = int(1000250001)
    structure_type_framebuffer_mixed_samples_combination_nv = int(1000250002)
    structure_type_physical_device_fragment_shader_interlock_features_ext = int(1000251000)
    structure_type_physical_device_ycbcr_image_arrays_features_ext = int(1000252000)
    structure_type_physical_device_provoking_vertex_features_ext = int(1000254000)
    structure_type_pipeline_rasterization_provoking_vertex_state_create_info_ext = int(1000254001)
    structure_type_physical_device_provoking_vertex_properties_ext = int(1000254002)
    structure_type_surface_full_screen_exclusive_info_ext = int(1000255000)
    structure_type_surface_capabilities_full_screen_exclusive_ext = int(1000255002)
    structure_type_surface_full_screen_exclusive_win32_info_ext = int(1000255001)
    structure_type_headless_surface_create_info_ext = int(1000256000)
    structure_type_physical_device_line_rasterization_features_ext = int(1000259000)
    structure_type_pipeline_rasterization_line_state_create_info_ext = int(1000259001)
    structure_type_physical_device_line_rasterization_properties_ext = int(1000259002)
    structure_type_physical_device_shader_atomic_float_features_ext = int(1000260000)
    structure_type_physical_device_index_type_uint8_features_ext = int(1000265000)
    structure_type_physical_device_extended_dynamic_state_features_ext = int(1000267000)
    structure_type_physical_device_pipeline_executable_properties_features_khr = int(1000269000)
    structure_type_pipeline_info_khr = int(1000269001)
    structure_type_pipeline_executable_properties_khr = int(1000269002)
    structure_type_pipeline_executable_info_khr = int(1000269003)
    structure_type_pipeline_executable_statistic_khr = int(1000269004)
    structure_type_pipeline_executable_internal_representation_khr = int(1000269005)
    structure_type_physical_device_host_image_copy_features_ext = int(1000270000)
    structure_type_physical_device_host_image_copy_properties_ext = int(1000270001)
    structure_type_memory_to_image_copy_ext = int(1000270002)
    structure_type_image_to_memory_copy_ext = int(1000270003)
    structure_type_copy_image_to_memory_info_ext = int(1000270004)
    structure_type_copy_memory_to_image_info_ext = int(1000270005)
    structure_type_host_image_layout_transition_info_ext = int(1000270006)
    structure_type_copy_image_to_image_info_ext = int(1000270007)
    structure_type_subresource_host_memcpy_size_ext = int(1000270008)
    structure_type_host_image_copy_device_performance_query_ext = int(1000270009)
    structure_type_memory_map_info_khr = int(1000271000)
    structure_type_memory_unmap_info_khr = int(1000271001)
    structure_type_physical_device_shader_atomic_float_2_features_ext = int(1000273000)
    structure_type_surface_present_mode_ext = int(1000274000)
    structure_type_surface_present_scaling_capabilities_ext = int(1000274001)
    structure_type_surface_present_mode_compatibility_ext = int(1000274002)
    structure_type_physical_device_swapchain_maintenance_1_features_ext = int(1000275000)
    structure_type_swapchain_present_fence_info_ext = int(1000275001)
    structure_type_swapchain_present_modes_create_info_ext = int(1000275002)
    structure_type_swapchain_present_mode_info_ext = int(1000275003)
    structure_type_swapchain_present_scaling_create_info_ext = int(1000275004)
    structure_type_release_swapchain_images_info_ext = int(1000275005)
    structure_type_physical_device_device_generated_commands_properties_nv = int(1000277000)
    structure_type_graphics_shader_group_create_info_nv = int(1000277001)
    structure_type_graphics_pipeline_shader_groups_create_info_nv = int(1000277002)
    structure_type_indirect_commands_layout_token_nv = int(1000277003)
    structure_type_indirect_commands_layout_create_info_nv = int(1000277004)
    structure_type_generated_commands_info_nv = int(1000277005)
    structure_type_generated_commands_memory_requirements_info_nv = int(1000277006)
    structure_type_physical_device_device_generated_commands_features_nv = int(1000277007)
    structure_type_physical_device_inherited_viewport_scissor_features_nv = int(1000278000)
    structure_type_command_buffer_inheritance_viewport_scissor_info_nv = int(1000278001)
    structure_type_physical_device_texel_buffer_alignment_features_ext = int(1000281000)
    structure_type_command_buffer_inheritance_render_pass_transform_info_qcom = int(1000282000)
    structure_type_render_pass_transform_begin_info_qcom = int(1000282001)
    structure_type_physical_device_depth_bias_control_features_ext = int(1000283000)
    structure_type_depth_bias_info_ext = int(1000283001)
    structure_type_depth_bias_representation_info_ext = int(1000283002)
    structure_type_physical_device_device_memory_report_features_ext = int(1000284000)
    structure_type_device_device_memory_report_create_info_ext = int(1000284001)
    structure_type_device_memory_report_callback_data_ext = int(1000284002)
    structure_type_physical_device_robustness_2_features_ext = int(1000286000)
    structure_type_physical_device_robustness_2_properties_ext = int(1000286001)
    structure_type_sampler_custom_border_color_create_info_ext = int(1000287000)
    structure_type_physical_device_custom_border_color_properties_ext = int(1000287001)
    structure_type_physical_device_custom_border_color_features_ext = int(1000287002)
    structure_type_pipeline_library_create_info_khr = int(1000290000)
    structure_type_physical_device_present_barrier_features_nv = int(1000292000)
    structure_type_surface_capabilities_present_barrier_nv = int(1000292001)
    structure_type_swapchain_present_barrier_create_info_nv = int(1000292002)
    structure_type_present_id_khr = int(1000294000)
    structure_type_physical_device_present_id_features_khr = int(1000294001)
    structure_type_physical_device_diagnostics_config_features_nv = int(1000300000)
    structure_type_device_diagnostics_config_create_info_nv = int(1000300001)
    structure_type_cuda_module_create_info_nv = int(1000307000)
    structure_type_cuda_function_create_info_nv = int(1000307001)
    structure_type_cuda_launch_info_nv = int(1000307002)
    structure_type_physical_device_cuda_kernel_launch_features_nv = int(1000307003)
    structure_type_physical_device_cuda_kernel_launch_properties_nv = int(1000307004)
    structure_type_query_low_latency_support_nv = int(1000310000)
    structure_type_export_metal_object_create_info_ext = int(1000311000)
    structure_type_export_metal_objects_info_ext = int(1000311001)
    structure_type_export_metal_device_info_ext = int(1000311002)
    structure_type_export_metal_command_queue_info_ext = int(1000311003)
    structure_type_export_metal_buffer_info_ext = int(1000311004)
    structure_type_import_metal_buffer_info_ext = int(1000311005)
    structure_type_export_metal_texture_info_ext = int(1000311006)
    structure_type_import_metal_texture_info_ext = int(1000311007)
    structure_type_export_metal_io_surface_info_ext = int(1000311008)
    structure_type_import_metal_io_surface_info_ext = int(1000311009)
    structure_type_export_metal_shared_event_info_ext = int(1000311010)
    structure_type_import_metal_shared_event_info_ext = int(1000311011)
    structure_type_queue_family_checkpoint_properties_2_nv = int(1000314008)
    structure_type_checkpoint_data_2_nv = int(1000314009)
    structure_type_physical_device_descriptor_buffer_properties_ext = int(1000316000)
    structure_type_physical_device_descriptor_buffer_density_map_properties_ext = int(1000316001)
    structure_type_physical_device_descriptor_buffer_features_ext = int(1000316002)
    structure_type_descriptor_address_info_ext = int(1000316003)
    structure_type_descriptor_get_info_ext = int(1000316004)
    structure_type_buffer_capture_descriptor_data_info_ext = int(1000316005)
    structure_type_image_capture_descriptor_data_info_ext = int(1000316006)
    structure_type_image_view_capture_descriptor_data_info_ext = int(1000316007)
    structure_type_sampler_capture_descriptor_data_info_ext = int(1000316008)
    structure_type_opaque_capture_descriptor_data_create_info_ext = int(1000316010)
    structure_type_descriptor_buffer_binding_info_ext = int(1000316011)
    structure_type_descriptor_buffer_binding_push_descriptor_buffer_handle_ext = int(1000316012)
    structure_type_acceleration_structure_capture_descriptor_data_info_ext = int(1000316009)
    structure_type_physical_device_graphics_pipeline_library_features_ext = int(1000320000)
    structure_type_physical_device_graphics_pipeline_library_properties_ext = int(1000320001)
    structure_type_graphics_pipeline_library_create_info_ext = int(1000320002)
    structure_type_physical_device_shader_early_and_late_fragment_tests_features_amd = int(1000321000)
    structure_type_physical_device_fragment_shader_barycentric_features_khr = int(1000203000)
    structure_type_physical_device_fragment_shader_barycentric_properties_khr = int(1000322000)
    structure_type_physical_device_shader_subgroup_uniform_control_flow_features_khr = int(1000323000)
    structure_type_physical_device_fragment_shading_rate_enums_properties_nv = int(1000326000)
    structure_type_physical_device_fragment_shading_rate_enums_features_nv = int(1000326001)
    structure_type_pipeline_fragment_shading_rate_enum_state_create_info_nv = int(1000326002)
    structure_type_acceleration_structure_geometry_motion_triangles_data_nv = int(1000327000)
    structure_type_physical_device_ray_tracing_motion_blur_features_nv = int(1000327001)
    structure_type_acceleration_structure_motion_info_nv = int(1000327002)
    structure_type_physical_device_mesh_shader_features_ext = int(1000328000)
    structure_type_physical_device_mesh_shader_properties_ext = int(1000328001)
    structure_type_physical_device_ycbcr_2_plane_444_formats_features_ext = int(1000330000)
    structure_type_physical_device_fragment_density_map_2_features_ext = int(1000332000)
    structure_type_physical_device_fragment_density_map_2_properties_ext = int(1000332001)
    structure_type_copy_command_transform_info_qcom = int(1000333000)
    structure_type_physical_device_workgroup_memory_explicit_layout_features_khr = int(1000336000)
    structure_type_physical_device_image_compression_control_features_ext = int(1000338000)
    structure_type_image_compression_control_ext = int(1000338001)
    structure_type_image_compression_properties_ext = int(1000338004)
    structure_type_physical_device_attachment_feedback_loop_layout_features_ext = int(1000339000)
    structure_type_physical_device_4444_formats_features_ext = int(1000340000)
    structure_type_physical_device_fault_features_ext = int(1000341000)
    structure_type_device_fault_counts_ext = int(1000341001)
    structure_type_device_fault_info_ext = int(1000341002)
    structure_type_physical_device_rgba10x6_formats_features_ext = int(1000344000)
    structure_type_directfb_surface_create_info_ext = int(1000346000)
    structure_type_physical_device_vertex_input_dynamic_state_features_ext = int(1000352000)
    structure_type_vertex_input_binding_description_2_ext = int(1000352001)
    structure_type_vertex_input_attribute_description_2_ext = int(1000352002)
    structure_type_physical_device_drm_properties_ext = int(1000353000)
    structure_type_physical_device_address_binding_report_features_ext = int(1000354000)
    structure_type_device_address_binding_callback_data_ext = int(1000354001)
    structure_type_physical_device_depth_clip_control_features_ext = int(1000355000)
    structure_type_pipeline_viewport_depth_clip_control_create_info_ext = int(1000355001)
    structure_type_physical_device_primitive_topology_list_restart_features_ext = int(1000356000)
    structure_type_import_memory_zircon_handle_info_fuchsia = int(1000364000)
    structure_type_memory_zircon_handle_properties_fuchsia = int(1000364001)
    structure_type_memory_get_zircon_handle_info_fuchsia = int(1000364002)
    structure_type_import_semaphore_zircon_handle_info_fuchsia = int(1000365000)
    structure_type_semaphore_get_zircon_handle_info_fuchsia = int(1000365001)
    structure_type_buffer_collection_create_info_fuchsia = int(1000366000)
    structure_type_import_memory_buffer_collection_fuchsia = int(1000366001)
    structure_type_buffer_collection_image_create_info_fuchsia = int(1000366002)
    structure_type_buffer_collection_properties_fuchsia = int(1000366003)
    structure_type_buffer_constraints_info_fuchsia = int(1000366004)
    structure_type_buffer_collection_buffer_create_info_fuchsia = int(1000366005)
    structure_type_image_constraints_info_fuchsia = int(1000366006)
    structure_type_image_format_constraints_info_fuchsia = int(1000366007)
    structure_type_sysmem_color_space_fuchsia = int(1000366008)
    structure_type_buffer_collection_constraints_info_fuchsia = int(1000366009)
    structure_type_subpass_shading_pipeline_create_info_huawei = int(1000369000)
    structure_type_physical_device_subpass_shading_features_huawei = int(1000369001)
    structure_type_physical_device_subpass_shading_properties_huawei = int(1000369002)
    structure_type_physical_device_invocation_mask_features_huawei = int(1000370000)
    structure_type_memory_get_remote_address_info_nv = int(1000371000)
    structure_type_physical_device_external_memory_rdma_features_nv = int(1000371001)
    structure_type_pipeline_properties_identifier_ext = int(1000372000)
    structure_type_physical_device_pipeline_properties_features_ext = int(1000372001)
    structure_type_physical_device_frame_boundary_features_ext = int(1000375000)
    structure_type_frame_boundary_ext = int(1000375001)
    structure_type_physical_device_multisampled_render_to_single_sampled_features_ext = int(1000376000)
    structure_type_subpass_resolve_performance_query_ext = int(1000376001)
    structure_type_multisampled_render_to_single_sampled_info_ext = int(1000376002)
    structure_type_physical_device_extended_dynamic_state_2_features_ext = int(1000377000)
    structure_type_screen_surface_create_info_qnx = int(1000378000)
    structure_type_physical_device_color_write_enable_features_ext = int(1000381000)
    structure_type_pipeline_color_write_create_info_ext = int(1000381001)
    structure_type_physical_device_primitives_generated_query_features_ext = int(1000382000)
    structure_type_physical_device_ray_tracing_maintenance_1_features_khr = int(1000386000)
    structure_type_physical_device_image_view_min_lod_features_ext = int(1000391000)
    structure_type_image_view_min_lod_create_info_ext = int(1000391001)
    structure_type_physical_device_multi_draw_features_ext = int(1000392000)
    structure_type_physical_device_multi_draw_properties_ext = int(1000392001)
    structure_type_physical_device_image_2d_view_of_3d_features_ext = int(1000393000)
    structure_type_physical_device_shader_tile_image_features_ext = int(1000395000)
    structure_type_physical_device_shader_tile_image_properties_ext = int(1000395001)
    structure_type_micromap_build_info_ext = int(1000396000)
    structure_type_micromap_version_info_ext = int(1000396001)
    structure_type_copy_micromap_info_ext = int(1000396002)
    structure_type_copy_micromap_to_memory_info_ext = int(1000396003)
    structure_type_copy_memory_to_micromap_info_ext = int(1000396004)
    structure_type_physical_device_opacity_micromap_features_ext = int(1000396005)
    structure_type_physical_device_opacity_micromap_properties_ext = int(1000396006)
    structure_type_micromap_create_info_ext = int(1000396007)
    structure_type_micromap_build_sizes_info_ext = int(1000396008)
    structure_type_acceleration_structure_triangles_opacity_micromap_ext = int(1000396009)
    structure_type_physical_device_cluster_culling_shader_features_huawei = int(1000404000)
    structure_type_physical_device_cluster_culling_shader_properties_huawei = int(1000404001)
    structure_type_physical_device_cluster_culling_shader_vrs_features_huawei = int(1000404002)
    structure_type_physical_device_border_color_swizzle_features_ext = int(1000411000)
    structure_type_sampler_border_color_component_mapping_create_info_ext = int(1000411001)
    structure_type_physical_device_pageable_device_local_memory_features_ext = int(1000412000)
    structure_type_physical_device_shader_core_properties_arm = int(1000415000)
    structure_type_device_queue_shader_core_control_create_info_arm = int(1000417000)
    structure_type_physical_device_scheduling_controls_features_arm = int(1000417001)
    structure_type_physical_device_scheduling_controls_properties_arm = int(1000417002)
    structure_type_physical_device_image_sliced_view_of_3d_features_ext = int(1000418000)
    structure_type_image_view_sliced_create_info_ext = int(1000418001)
    structure_type_physical_device_descriptor_set_host_mapping_features_valve = int(1000420000)
    structure_type_descriptor_set_binding_reference_valve = int(1000420001)
    structure_type_descriptor_set_layout_host_mapping_info_valve = int(1000420002)
    structure_type_physical_device_depth_clamp_zero_one_features_ext = int(1000421000)
    structure_type_physical_device_non_seamless_cube_map_features_ext = int(1000422000)
    structure_type_physical_device_render_pass_striped_features_arm = int(1000424000)
    structure_type_physical_device_render_pass_striped_properties_arm = int(1000424001)
    structure_type_render_pass_stripe_begin_info_arm = int(1000424002)
    structure_type_render_pass_stripe_info_arm = int(1000424003)
    structure_type_render_pass_stripe_submit_info_arm = int(1000424004)
    structure_type_physical_device_fragment_density_map_offset_features_qcom = int(1000425000)
    structure_type_physical_device_fragment_density_map_offset_properties_qcom = int(1000425001)
    structure_type_subpass_fragment_density_map_offset_end_info_qcom = int(1000425002)
    structure_type_physical_device_copy_memory_indirect_features_nv = int(1000426000)
    structure_type_physical_device_copy_memory_indirect_properties_nv = int(1000426001)
    structure_type_physical_device_memory_decompression_features_nv = int(1000427000)
    structure_type_physical_device_memory_decompression_properties_nv = int(1000427001)
    structure_type_physical_device_device_generated_commands_compute_features_nv = int(1000428000)
    structure_type_compute_pipeline_indirect_buffer_info_nv = int(1000428001)
    structure_type_pipeline_indirect_device_address_info_nv = int(1000428002)
    structure_type_physical_device_linear_color_attachment_features_nv = int(1000430000)
    structure_type_physical_device_image_compression_control_swapchain_features_ext = int(1000437000)
    structure_type_physical_device_image_processing_features_qcom = int(1000440000)
    structure_type_physical_device_image_processing_properties_qcom = int(1000440001)
    structure_type_image_view_sample_weight_create_info_qcom = int(1000440002)
    structure_type_physical_device_nested_command_buffer_features_ext = int(1000451000)
    structure_type_physical_device_nested_command_buffer_properties_ext = int(1000451001)
    structure_type_external_memory_acquire_unmodified_ext = int(1000453000)
    structure_type_physical_device_extended_dynamic_state_3_features_ext = int(1000455000)
    structure_type_physical_device_extended_dynamic_state_3_properties_ext = int(1000455001)
    structure_type_physical_device_subpass_merge_feedback_features_ext = int(1000458000)
    structure_type_render_pass_creation_control_ext = int(1000458001)
    structure_type_render_pass_creation_feedback_create_info_ext = int(1000458002)
    structure_type_render_pass_subpass_feedback_create_info_ext = int(1000458003)
    structure_type_direct_driver_loading_info_lunarg = int(1000459000)
    structure_type_direct_driver_loading_list_lunarg = int(1000459001)
    structure_type_physical_device_shader_module_identifier_features_ext = int(1000462000)
    structure_type_physical_device_shader_module_identifier_properties_ext = int(1000462001)
    structure_type_pipeline_shader_stage_module_identifier_create_info_ext = int(1000462002)
    structure_type_shader_module_identifier_ext = int(1000462003)
    structure_type_physical_device_rasterization_order_attachment_access_features_ext = int(1000342000)
    structure_type_physical_device_optical_flow_features_nv = int(1000464000)
    structure_type_physical_device_optical_flow_properties_nv = int(1000464001)
    structure_type_optical_flow_image_format_info_nv = int(1000464002)
    structure_type_optical_flow_image_format_properties_nv = int(1000464003)
    structure_type_optical_flow_session_create_info_nv = int(1000464004)
    structure_type_optical_flow_execute_info_nv = int(1000464005)
    structure_type_optical_flow_session_create_private_data_info_nv = int(1000464010)
    structure_type_physical_device_legacy_dithering_features_ext = int(1000465000)
    structure_type_physical_device_pipeline_protected_access_features_ext = int(1000466000)
    structure_type_physical_device_external_format_resolve_features_android = int(1000468000)
    structure_type_physical_device_external_format_resolve_properties_android = int(1000468001)
    structure_type_android_hardware_buffer_format_resolve_properties_android = int(1000468002)
    structure_type_physical_device_maintenance_5_features_khr = int(1000470000)
    structure_type_physical_device_maintenance_5_properties_khr = int(1000470001)
    structure_type_rendering_area_info_khr = int(1000470003)
    structure_type_device_image_subresource_info_khr = int(1000470004)
    structure_type_subresource_layout_2_khr = int(1000338002)
    structure_type_image_subresource_2_khr = int(1000338003)
    structure_type_pipeline_create_flags_2_create_info_khr = int(1000470005)
    structure_type_buffer_usage_flags_2_create_info_khr = int(1000470006)
    structure_type_physical_device_ray_tracing_position_fetch_features_khr = int(1000481000)
    structure_type_physical_device_shader_object_features_ext = int(1000482000)
    structure_type_physical_device_shader_object_properties_ext = int(1000482001)
    structure_type_shader_create_info_ext = int(1000482002)
    structure_type_physical_device_tile_properties_features_qcom = int(1000484000)
    structure_type_tile_properties_qcom = int(1000484001)
    structure_type_physical_device_amigo_profiling_features_sec = int(1000485000)
    structure_type_amigo_profiling_submit_info_sec = int(1000485001)
    structure_type_physical_device_multiview_per_view_viewports_features_qcom = int(1000488000)
    structure_type_physical_device_ray_tracing_invocation_reorder_features_nv = int(1000490000)
    structure_type_physical_device_ray_tracing_invocation_reorder_properties_nv = int(1000490001)
    structure_type_physical_device_extended_sparse_address_space_features_nv = int(1000492000)
    structure_type_physical_device_extended_sparse_address_space_properties_nv = int(1000492001)
    structure_type_physical_device_mutable_descriptor_type_features_ext = int(1000351000)
    structure_type_mutable_descriptor_type_create_info_ext = int(1000351002)
    structure_type_layer_settings_create_info_ext = int(1000496000)
    structure_type_physical_device_shader_core_builtins_features_arm = int(1000497000)
    structure_type_physical_device_shader_core_builtins_properties_arm = int(1000497001)
    structure_type_physical_device_pipeline_library_group_handles_features_ext = int(1000498000)
    structure_type_physical_device_dynamic_rendering_unused_attachments_features_ext = int(1000499000)
    structure_type_latency_sleep_mode_info_nv = int(1000505000)
    structure_type_latency_sleep_info_nv = int(1000505001)
    structure_type_set_latency_marker_info_nv = int(1000505002)
    structure_type_get_latency_marker_info_nv = int(1000505003)
    structure_type_latency_timings_frame_report_nv = int(1000505004)
    structure_type_latency_submission_present_id_nv = int(1000505005)
    structure_type_out_of_band_queue_type_info_nv = int(1000505006)
    structure_type_swapchain_latency_create_info_nv = int(1000505007)
    structure_type_latency_surface_capabilities_nv = int(1000505008)
    structure_type_physical_device_cooperative_matrix_features_khr = int(1000506000)
    structure_type_cooperative_matrix_properties_khr = int(1000506001)
    structure_type_physical_device_cooperative_matrix_properties_khr = int(1000506002)
    structure_type_physical_device_multiview_per_view_render_areas_features_qcom = int(1000510000)
    structure_type_multiview_per_view_render_areas_render_pass_begin_info_qcom = int(1000510001)
    structure_type_physical_device_image_processing_2_features_qcom = int(1000518000)
    structure_type_physical_device_image_processing_2_properties_qcom = int(1000518001)
    structure_type_sampler_block_match_window_create_info_qcom = int(1000518002)
    structure_type_sampler_cubic_weights_create_info_qcom = int(1000519000)
    structure_type_physical_device_cubic_weights_features_qcom = int(1000519001)
    structure_type_blit_image_cubic_weights_info_qcom = int(1000519002)
    structure_type_physical_device_ycbcr_degamma_features_qcom = int(1000520000)
    structure_type_sampler_ycbcr_conversion_ycbcr_degamma_create_info_qcom = int(1000520001)
    structure_type_physical_device_cubic_clamp_features_qcom = int(1000521000)
    structure_type_physical_device_attachment_feedback_loop_dynamic_state_features_ext = int(1000524000)
    structure_type_screen_buffer_properties_qnx = int(1000529000)
    structure_type_screen_buffer_format_properties_qnx = int(1000529001)
    structure_type_import_screen_buffer_info_qnx = int(1000529002)
    structure_type_external_format_qnx = int(1000529003)
    structure_type_physical_device_external_memory_screen_buffer_features_qnx = int(1000529004)
    structure_type_physical_device_layered_driver_properties_msft = int(1000530000)
    structure_type_physical_device_descriptor_pool_overallocation_features_nv = int(1000546000)
    structure_type_max_enum = int(0x7FFFFFFF)
}


pub enum PipelineCacheHeaderVersion {
    pipeline_cache_header_version_one = int(1)
    pipeline_cache_header_version_max_enum = int(0x7FFFFFFF)
}


pub enum ImageLayout {
    image_layout_undefined = int(0)
    image_layout_general = int(1)
    image_layout_color_attachment_optimal = int(2)
    image_layout_depth_stencil_attachment_optimal = int(3)
    image_layout_depth_stencil_read_only_optimal = int(4)
    image_layout_shader_read_only_optimal = int(5)
    image_layout_transfer_src_optimal = int(6)
    image_layout_transfer_dst_optimal = int(7)
    image_layout_preinitialized = int(8)
    image_layout_depth_read_only_stencil_attachment_optimal = int(1000117000)
    image_layout_depth_attachment_stencil_read_only_optimal = int(1000117001)
    image_layout_depth_attachment_optimal = int(1000241000)
    image_layout_depth_read_only_optimal = int(1000241001)
    image_layout_stencil_attachment_optimal = int(1000241002)
    image_layout_stencil_read_only_optimal = int(1000241003)
    image_layout_read_only_optimal = int(1000314000)
    image_layout_attachment_optimal = int(1000314001)
    image_layout_present_src_khr = int(1000001002)
    image_layout_video_decode_dst_khr = int(1000024000)
    image_layout_video_decode_src_khr = int(1000024001)
    image_layout_video_decode_dpb_khr = int(1000024002)
    image_layout_shared_present_khr = int(1000111000)
    image_layout_fragment_density_map_optimal_ext = int(1000218000)
    image_layout_fragment_shading_rate_attachment_optimal_khr = int(1000164003)
    image_layout_attachment_feedback_loop_optimal_ext = int(1000339000)
    image_layout_max_enum = int(0x7FFFFFFF)
}


pub enum ObjectType {
    object_type_unknown = int(0)
    object_type_instance = int(1)
    object_type_physical_device = int(2)
    object_type_device = int(3)
    object_type_queue = int(4)
    object_type_semaphore = int(5)
    object_type_command_buffer = int(6)
    object_type_fence = int(7)
    object_type_device_memory = int(8)
    object_type_buffer = int(9)
    object_type_image = int(10)
    object_type_event = int(11)
    object_type_query_pool = int(12)
    object_type_buffer_view = int(13)
    object_type_image_view = int(14)
    object_type_shader_module = int(15)
    object_type_pipeline_cache = int(16)
    object_type_pipeline_layout = int(17)
    object_type_render_pass = int(18)
    object_type_pipeline = int(19)
    object_type_descriptor_set_layout = int(20)
    object_type_sampler = int(21)
    object_type_descriptor_pool = int(22)
    object_type_descriptor_set = int(23)
    object_type_framebuffer = int(24)
    object_type_command_pool = int(25)
    object_type_sampler_ycbcr_conversion = int(1000156000)
    object_type_descriptor_update_template = int(1000085000)
    object_type_private_data_slot = int(1000295000)
    object_type_surface_khr = int(1000000000)
    object_type_swapchain_khr = int(1000001000)
    object_type_display_khr = int(1000002000)
    object_type_display_mode_khr = int(1000002001)
    object_type_debug_report_callback_ext = int(1000011000)
    object_type_video_session_khr = int(1000023000)
    object_type_video_session_parameters_khr = int(1000023001)
    object_type_cu_module_nvx = int(1000029000)
    object_type_cu_function_nvx = int(1000029001)
    object_type_debug_utils_messenger_ext = int(1000128000)
    object_type_acceleration_structure_khr = int(1000150000)
    object_type_validation_cache_ext = int(1000160000)
    object_type_acceleration_structure_nv = int(1000165000)
    object_type_performance_configuration_intel = int(1000210000)
    object_type_deferred_operation_khr = int(1000268000)
    object_type_indirect_commands_layout_nv = int(1000277000)
    object_type_cuda_module_nv = int(1000307000)
    object_type_cuda_function_nv = int(1000307001)
    object_type_buffer_collection_fuchsia = int(1000366000)
    object_type_micromap_ext = int(1000396000)
    object_type_optical_flow_session_nv = int(1000464000)
    object_type_shader_ext = int(1000482000)
    object_type_max_enum = int(0x7FFFFFFF)
}


pub enum VendorId {
    vendor_id_viv = int(0x10001)
    vendor_id_vsi = int(0x10002)
    vendor_id_kazan = int(0x10003)
    vendor_id_codeplay = int(0x10004)
    vendor_id_mesa = int(0x10005)
    vendor_id_pocl = int(0x10006)
    vendor_id_mobileye = int(0x10007)
    vendor_id_max_enum = int(0x7FFFFFFF)
}


pub enum SystemAllocationScope {
    system_allocation_scope_command = int(0)
    system_allocation_scope_object = int(1)
    system_allocation_scope_cache = int(2)
    system_allocation_scope_device = int(3)
    system_allocation_scope_instance = int(4)
    system_allocation_scope_max_enum = int(0x7FFFFFFF)
}


pub enum InternalAllocationType {
    internal_allocation_type_executable = int(0)
    internal_allocation_type_max_enum = int(0x7FFFFFFF)
}


pub enum Format {
    format_undefined = int(0)
    format_r4g4_unorm_pack8 = int(1)
    format_r4g4b4a4_unorm_pack16 = int(2)
    format_b4g4r4a4_unorm_pack16 = int(3)
    format_r5g6b5_unorm_pack16 = int(4)
    format_b5g6r5_unorm_pack16 = int(5)
    format_r5g5b5a1_unorm_pack16 = int(6)
    format_b5g5r5a1_unorm_pack16 = int(7)
    format_a1r5g5b5_unorm_pack16 = int(8)
    format_r8_unorm = int(9)
    format_r8_snorm = int(10)
    format_r8_uscaled = int(11)
    format_r8_sscaled = int(12)
    format_r8_uint = int(13)
    format_r8_sint = int(14)
    format_r8_srgb = int(15)
    format_r8g8_unorm = int(16)
    format_r8g8_snorm = int(17)
    format_r8g8_uscaled = int(18)
    format_r8g8_sscaled = int(19)
    format_r8g8_uint = int(20)
    format_r8g8_sint = int(21)
    format_r8g8_srgb = int(22)
    format_r8g8b8_unorm = int(23)
    format_r8g8b8_snorm = int(24)
    format_r8g8b8_uscaled = int(25)
    format_r8g8b8_sscaled = int(26)
    format_r8g8b8_uint = int(27)
    format_r8g8b8_sint = int(28)
    format_r8g8b8_srgb = int(29)
    format_b8g8r8_unorm = int(30)
    format_b8g8r8_snorm = int(31)
    format_b8g8r8_uscaled = int(32)
    format_b8g8r8_sscaled = int(33)
    format_b8g8r8_uint = int(34)
    format_b8g8r8_sint = int(35)
    format_b8g8r8_srgb = int(36)
    format_r8g8b8a8_unorm = int(37)
    format_r8g8b8a8_snorm = int(38)
    format_r8g8b8a8_uscaled = int(39)
    format_r8g8b8a8_sscaled = int(40)
    format_r8g8b8a8_uint = int(41)
    format_r8g8b8a8_sint = int(42)
    format_r8g8b8a8_srgb = int(43)
    format_b8g8r8a8_unorm = int(44)
    format_b8g8r8a8_snorm = int(45)
    format_b8g8r8a8_uscaled = int(46)
    format_b8g8r8a8_sscaled = int(47)
    format_b8g8r8a8_uint = int(48)
    format_b8g8r8a8_sint = int(49)
    format_b8g8r8a8_srgb = int(50)
    format_a8b8g8r8_unorm_pack32 = int(51)
    format_a8b8g8r8_snorm_pack32 = int(52)
    format_a8b8g8r8_uscaled_pack32 = int(53)
    format_a8b8g8r8_sscaled_pack32 = int(54)
    format_a8b8g8r8_uint_pack32 = int(55)
    format_a8b8g8r8_sint_pack32 = int(56)
    format_a8b8g8r8_srgb_pack32 = int(57)
    format_a2r10g10b10_unorm_pack32 = int(58)
    format_a2r10g10b10_snorm_pack32 = int(59)
    format_a2r10g10b10_uscaled_pack32 = int(60)
    format_a2r10g10b10_sscaled_pack32 = int(61)
    format_a2r10g10b10_uint_pack32 = int(62)
    format_a2r10g10b10_sint_pack32 = int(63)
    format_a2b10g10r10_unorm_pack32 = int(64)
    format_a2b10g10r10_snorm_pack32 = int(65)
    format_a2b10g10r10_uscaled_pack32 = int(66)
    format_a2b10g10r10_sscaled_pack32 = int(67)
    format_a2b10g10r10_uint_pack32 = int(68)
    format_a2b10g10r10_sint_pack32 = int(69)
    format_r16_unorm = int(70)
    format_r16_snorm = int(71)
    format_r16_uscaled = int(72)
    format_r16_sscaled = int(73)
    format_r16_uint = int(74)
    format_r16_sint = int(75)
    format_r16_sfloat = int(76)
    format_r16g16_unorm = int(77)
    format_r16g16_snorm = int(78)
    format_r16g16_uscaled = int(79)
    format_r16g16_sscaled = int(80)
    format_r16g16_uint = int(81)
    format_r16g16_sint = int(82)
    format_r16g16_sfloat = int(83)
    format_r16g16b16_unorm = int(84)
    format_r16g16b16_snorm = int(85)
    format_r16g16b16_uscaled = int(86)
    format_r16g16b16_sscaled = int(87)
    format_r16g16b16_uint = int(88)
    format_r16g16b16_sint = int(89)
    format_r16g16b16_sfloat = int(90)
    format_r16g16b16a16_unorm = int(91)
    format_r16g16b16a16_snorm = int(92)
    format_r16g16b16a16_uscaled = int(93)
    format_r16g16b16a16_sscaled = int(94)
    format_r16g16b16a16_uint = int(95)
    format_r16g16b16a16_sint = int(96)
    format_r16g16b16a16_sfloat = int(97)
    format_r32_uint = int(98)
    format_r32_sint = int(99)
    format_r32_sfloat = int(100)
    format_r32g32_uint = int(101)
    format_r32g32_sint = int(102)
    format_r32g32_sfloat = int(103)
    format_r32g32b32_uint = int(104)
    format_r32g32b32_sint = int(105)
    format_r32g32b32_sfloat = int(106)
    format_r32g32b32a32_uint = int(107)
    format_r32g32b32a32_sint = int(108)
    format_r32g32b32a32_sfloat = int(109)
    format_r64_uint = int(110)
    format_r64_sint = int(111)
    format_r64_sfloat = int(112)
    format_r64g64_uint = int(113)
    format_r64g64_sint = int(114)
    format_r64g64_sfloat = int(115)
    format_r64g64b64_uint = int(116)
    format_r64g64b64_sint = int(117)
    format_r64g64b64_sfloat = int(118)
    format_r64g64b64a64_uint = int(119)
    format_r64g64b64a64_sint = int(120)
    format_r64g64b64a64_sfloat = int(121)
    format_b10g11r11_ufloat_pack32 = int(122)
    format_e5b9g9r9_ufloat_pack32 = int(123)
    format_d16_unorm = int(124)
    format_x8_d24_unorm_pack32 = int(125)
    format_d32_sfloat = int(126)
    format_s8_uint = int(127)
    format_d16_unorm_s8_uint = int(128)
    format_d24_unorm_s8_uint = int(129)
    format_d32_sfloat_s8_uint = int(130)
    format_bc1_rgb_unorm_block = int(131)
    format_bc1_rgb_srgb_block = int(132)
    format_bc1_rgba_unorm_block = int(133)
    format_bc1_rgba_srgb_block = int(134)
    format_bc2_unorm_block = int(135)
    format_bc2_srgb_block = int(136)
    format_bc3_unorm_block = int(137)
    format_bc3_srgb_block = int(138)
    format_bc4_unorm_block = int(139)
    format_bc4_snorm_block = int(140)
    format_bc5_unorm_block = int(141)
    format_bc5_snorm_block = int(142)
    format_bc6h_ufloat_block = int(143)
    format_bc6h_sfloat_block = int(144)
    format_bc7_unorm_block = int(145)
    format_bc7_srgb_block = int(146)
    format_etc2_r8g8b8_unorm_block = int(147)
    format_etc2_r8g8b8_srgb_block = int(148)
    format_etc2_r8g8b8a1_unorm_block = int(149)
    format_etc2_r8g8b8a1_srgb_block = int(150)
    format_etc2_r8g8b8a8_unorm_block = int(151)
    format_etc2_r8g8b8a8_srgb_block = int(152)
    format_eac_r11_unorm_block = int(153)
    format_eac_r11_snorm_block = int(154)
    format_eac_r11g11_unorm_block = int(155)
    format_eac_r11g11_snorm_block = int(156)
    format_astc_4x4_unorm_block = int(157)
    format_astc_4x4_srgb_block = int(158)
    format_astc_5x4_unorm_block = int(159)
    format_astc_5x4_srgb_block = int(160)
    format_astc_5x5_unorm_block = int(161)
    format_astc_5x5_srgb_block = int(162)
    format_astc_6x5_unorm_block = int(163)
    format_astc_6x5_srgb_block = int(164)
    format_astc_6x6_unorm_block = int(165)
    format_astc_6x6_srgb_block = int(166)
    format_astc_8x5_unorm_block = int(167)
    format_astc_8x5_srgb_block = int(168)
    format_astc_8x6_unorm_block = int(169)
    format_astc_8x6_srgb_block = int(170)
    format_astc_8x8_unorm_block = int(171)
    format_astc_8x8_srgb_block = int(172)
    format_astc_10x5_unorm_block = int(173)
    format_astc_10x5_srgb_block = int(174)
    format_astc_10x6_unorm_block = int(175)
    format_astc_10x6_srgb_block = int(176)
    format_astc_10x8_unorm_block = int(177)
    format_astc_10x8_srgb_block = int(178)
    format_astc_10x10_unorm_block = int(179)
    format_astc_10x10_srgb_block = int(180)
    format_astc_12x10_unorm_block = int(181)
    format_astc_12x10_srgb_block = int(182)
    format_astc_12x12_unorm_block = int(183)
    format_astc_12x12_srgb_block = int(184)
    format_g8b8g8r8_422_unorm = int(1000156000)
    format_b8g8r8g8_422_unorm = int(1000156001)
    format_g8_b8_r8_3plane_420_unorm = int(1000156002)
    format_g8_b8r8_2plane_420_unorm = int(1000156003)
    format_g8_b8_r8_3plane_422_unorm = int(1000156004)
    format_g8_b8r8_2plane_422_unorm = int(1000156005)
    format_g8_b8_r8_3plane_444_unorm = int(1000156006)
    format_r10x6_unorm_pack16 = int(1000156007)
    format_r10x6g10x6_unorm_2pack16 = int(1000156008)
    format_r10x6g10x6b10x6a10x6_unorm_4pack16 = int(1000156009)
    format_g10x6b10x6g10x6r10x6_422_unorm_4pack16 = int(1000156010)
    format_b10x6g10x6r10x6g10x6_422_unorm_4pack16 = int(1000156011)
    format_g10x6_b10x6_r10x6_3plane_420_unorm_3pack16 = int(1000156012)
    format_g10x6_b10x6r10x6_2plane_420_unorm_3pack16 = int(1000156013)
    format_g10x6_b10x6_r10x6_3plane_422_unorm_3pack16 = int(1000156014)
    format_g10x6_b10x6r10x6_2plane_422_unorm_3pack16 = int(1000156015)
    format_g10x6_b10x6_r10x6_3plane_444_unorm_3pack16 = int(1000156016)
    format_r12x4_unorm_pack16 = int(1000156017)
    format_r12x4g12x4_unorm_2pack16 = int(1000156018)
    format_r12x4g12x4b12x4a12x4_unorm_4pack16 = int(1000156019)
    format_g12x4b12x4g12x4r12x4_422_unorm_4pack16 = int(1000156020)
    format_b12x4g12x4r12x4g12x4_422_unorm_4pack16 = int(1000156021)
    format_g12x4_b12x4_r12x4_3plane_420_unorm_3pack16 = int(1000156022)
    format_g12x4_b12x4r12x4_2plane_420_unorm_3pack16 = int(1000156023)
    format_g12x4_b12x4_r12x4_3plane_422_unorm_3pack16 = int(1000156024)
    format_g12x4_b12x4r12x4_2plane_422_unorm_3pack16 = int(1000156025)
    format_g12x4_b12x4_r12x4_3plane_444_unorm_3pack16 = int(1000156026)
    format_g16b16g16r16_422_unorm = int(1000156027)
    format_b16g16r16g16_422_unorm = int(1000156028)
    format_g16_b16_r16_3plane_420_unorm = int(1000156029)
    format_g16_b16r16_2plane_420_unorm = int(1000156030)
    format_g16_b16_r16_3plane_422_unorm = int(1000156031)
    format_g16_b16r16_2plane_422_unorm = int(1000156032)
    format_g16_b16_r16_3plane_444_unorm = int(1000156033)
    format_g8_b8r8_2plane_444_unorm = int(1000330000)
    format_g10x6_b10x6r10x6_2plane_444_unorm_3pack16 = int(1000330001)
    format_g12x4_b12x4r12x4_2plane_444_unorm_3pack16 = int(1000330002)
    format_g16_b16r16_2plane_444_unorm = int(1000330003)
    format_a4r4g4b4_unorm_pack16 = int(1000340000)
    format_a4b4g4r4_unorm_pack16 = int(1000340001)
    format_astc_4x4_sfloat_block = int(1000066000)
    format_astc_5x4_sfloat_block = int(1000066001)
    format_astc_5x5_sfloat_block = int(1000066002)
    format_astc_6x5_sfloat_block = int(1000066003)
    format_astc_6x6_sfloat_block = int(1000066004)
    format_astc_8x5_sfloat_block = int(1000066005)
    format_astc_8x6_sfloat_block = int(1000066006)
    format_astc_8x8_sfloat_block = int(1000066007)
    format_astc_10x5_sfloat_block = int(1000066008)
    format_astc_10x6_sfloat_block = int(1000066009)
    format_astc_10x8_sfloat_block = int(1000066010)
    format_astc_10x10_sfloat_block = int(1000066011)
    format_astc_12x10_sfloat_block = int(1000066012)
    format_astc_12x12_sfloat_block = int(1000066013)
    format_pvrtc1_2bpp_unorm_block_img = int(1000054000)
    format_pvrtc1_4bpp_unorm_block_img = int(1000054001)
    format_pvrtc2_2bpp_unorm_block_img = int(1000054002)
    format_pvrtc2_4bpp_unorm_block_img = int(1000054003)
    format_pvrtc1_2bpp_srgb_block_img = int(1000054004)
    format_pvrtc1_4bpp_srgb_block_img = int(1000054005)
    format_pvrtc2_2bpp_srgb_block_img = int(1000054006)
    format_pvrtc2_4bpp_srgb_block_img = int(1000054007)
    format_r16g16_s10_5_nv = int(1000464000)
    format_a1b5g5r5_unorm_pack16_khr = int(1000470000)
    format_a8_unorm_khr = int(1000470001)
    format_max_enum = int(0x7FFFFFFF)
}


pub enum ImageTiling {
    image_tiling_optimal = int(0)
    image_tiling_linear = int(1)
    image_tiling_drm_format_modifier_ext = int(1000158000)
    image_tiling_max_enum = int(0x7FFFFFFF)
}


pub enum ImageType {
    image_type_1d = int(0)
    image_type_2d = int(1)
    image_type_3d = int(2)
    image_type_max_enum = int(0x7FFFFFFF)
}


pub enum PhysicalDeviceType {
    physical_device_type_other = int(0)
    physical_device_type_integrated_gpu = int(1)
    physical_device_type_discrete_gpu = int(2)
    physical_device_type_virtual_gpu = int(3)
    physical_device_type_cpu = int(4)
    physical_device_type_max_enum = int(0x7FFFFFFF)
}


pub enum QueryType {
    query_type_occlusion = int(0)
    query_type_pipeline_statistics = int(1)
    query_type_timestamp = int(2)
    query_type_result_status_only_khr = int(1000023000)
    query_type_transform_feedback_stream_ext = int(1000028004)
    query_type_performance_query_khr = int(1000116000)
    query_type_acceleration_structure_compacted_size_khr = int(1000150000)
    query_type_acceleration_structure_serialization_size_khr = int(1000150001)
    query_type_acceleration_structure_compacted_size_nv = int(1000165000)
    query_type_performance_query_intel = int(1000210000)
    query_type_mesh_primitives_generated_ext = int(1000328000)
    query_type_primitives_generated_ext = int(1000382000)
    query_type_acceleration_structure_serialization_bottom_level_pointers_khr = int(1000386000)
    query_type_acceleration_structure_size_khr = int(1000386001)
    query_type_micromap_serialization_size_ext = int(1000396000)
    query_type_micromap_compacted_size_ext = int(1000396001)
    query_type_max_enum = int(0x7FFFFFFF)
}


pub enum SharingMode {
    sharing_mode_exclusive = int(0)
    sharing_mode_concurrent = int(1)
    sharing_mode_max_enum = int(0x7FFFFFFF)
}


pub enum ComponentSwizzle {
    component_swizzle_identity = int(0)
    component_swizzle_zero = int(1)
    component_swizzle_one = int(2)
    component_swizzle_r = int(3)
    component_swizzle_g = int(4)
    component_swizzle_b = int(5)
    component_swizzle_a = int(6)
    component_swizzle_max_enum = int(0x7FFFFFFF)
}


pub enum ImageViewType {
    image_view_type_1d = int(0)
    image_view_type_2d = int(1)
    image_view_type_3d = int(2)
    image_view_type_cube = int(3)
    image_view_type_1d_array = int(4)
    image_view_type_2d_array = int(5)
    image_view_type_cube_array = int(6)
    image_view_type_max_enum = int(0x7FFFFFFF)
}


pub enum BlendFactor {
    blend_factor_zero = int(0)
    blend_factor_one = int(1)
    blend_factor_src_color = int(2)
    blend_factor_one_minus_src_color = int(3)
    blend_factor_dst_color = int(4)
    blend_factor_one_minus_dst_color = int(5)
    blend_factor_src_alpha = int(6)
    blend_factor_one_minus_src_alpha = int(7)
    blend_factor_dst_alpha = int(8)
    blend_factor_one_minus_dst_alpha = int(9)
    blend_factor_constant_color = int(10)
    blend_factor_one_minus_constant_color = int(11)
    blend_factor_constant_alpha = int(12)
    blend_factor_one_minus_constant_alpha = int(13)
    blend_factor_src_alpha_saturate = int(14)
    blend_factor_src1_color = int(15)
    blend_factor_one_minus_src1_color = int(16)
    blend_factor_src1_alpha = int(17)
    blend_factor_one_minus_src1_alpha = int(18)
    blend_factor_max_enum = int(0x7FFFFFFF)
}


pub enum BlendOp {
    blend_op_add = int(0)
    blend_op_subtract = int(1)
    blend_op_reverse_subtract = int(2)
    blend_op_min = int(3)
    blend_op_max = int(4)
    blend_op_zero_ext = int(1000148000)
    blend_op_src_ext = int(1000148001)
    blend_op_dst_ext = int(1000148002)
    blend_op_src_over_ext = int(1000148003)
    blend_op_dst_over_ext = int(1000148004)
    blend_op_src_in_ext = int(1000148005)
    blend_op_dst_in_ext = int(1000148006)
    blend_op_src_out_ext = int(1000148007)
    blend_op_dst_out_ext = int(1000148008)
    blend_op_src_atop_ext = int(1000148009)
    blend_op_dst_atop_ext = int(1000148010)
    blend_op_xor_ext = int(1000148011)
    blend_op_multiply_ext = int(1000148012)
    blend_op_screen_ext = int(1000148013)
    blend_op_overlay_ext = int(1000148014)
    blend_op_darken_ext = int(1000148015)
    blend_op_lighten_ext = int(1000148016)
    blend_op_colordodge_ext = int(1000148017)
    blend_op_colorburn_ext = int(1000148018)
    blend_op_hardlight_ext = int(1000148019)
    blend_op_softlight_ext = int(1000148020)
    blend_op_difference_ext = int(1000148021)
    blend_op_exclusion_ext = int(1000148022)
    blend_op_invert_ext = int(1000148023)
    blend_op_invert_rgb_ext = int(1000148024)
    blend_op_lineardodge_ext = int(1000148025)
    blend_op_linearburn_ext = int(1000148026)
    blend_op_vividlight_ext = int(1000148027)
    blend_op_linearlight_ext = int(1000148028)
    blend_op_pinlight_ext = int(1000148029)
    blend_op_hardmix_ext = int(1000148030)
    blend_op_hsl_hue_ext = int(1000148031)
    blend_op_hsl_saturation_ext = int(1000148032)
    blend_op_hsl_color_ext = int(1000148033)
    blend_op_hsl_luminosity_ext = int(1000148034)
    blend_op_plus_ext = int(1000148035)
    blend_op_plus_clamped_ext = int(1000148036)
    blend_op_plus_clamped_alpha_ext = int(1000148037)
    blend_op_plus_darker_ext = int(1000148038)
    blend_op_minus_ext = int(1000148039)
    blend_op_minus_clamped_ext = int(1000148040)
    blend_op_contrast_ext = int(1000148041)
    blend_op_invert_ovg_ext = int(1000148042)
    blend_op_red_ext = int(1000148043)
    blend_op_green_ext = int(1000148044)
    blend_op_blue_ext = int(1000148045)
    blend_op_max_enum = int(0x7FFFFFFF)
}


pub enum CompareOp {
    compare_op_never = int(0)
    compare_op_less = int(1)
    compare_op_equal = int(2)
    compare_op_less_or_equal = int(3)
    compare_op_greater = int(4)
    compare_op_not_equal = int(5)
    compare_op_greater_or_equal = int(6)
    compare_op_always = int(7)
    compare_op_max_enum = int(0x7FFFFFFF)
}


pub enum DynamicState {
    dynamic_state_viewport = int(0)
    dynamic_state_scissor = int(1)
    dynamic_state_line_width = int(2)
    dynamic_state_depth_bias = int(3)
    dynamic_state_blend_constants = int(4)
    dynamic_state_depth_bounds = int(5)
    dynamic_state_stencil_compare_mask = int(6)
    dynamic_state_stencil_write_mask = int(7)
    dynamic_state_stencil_reference = int(8)
    dynamic_state_cull_mode = int(1000267000)
    dynamic_state_front_face = int(1000267001)
    dynamic_state_primitive_topology = int(1000267002)
    dynamic_state_viewport_with_count = int(1000267003)
    dynamic_state_scissor_with_count = int(1000267004)
    dynamic_state_vertex_input_binding_stride = int(1000267005)
    dynamic_state_depth_test_enable = int(1000267006)
    dynamic_state_depth_write_enable = int(1000267007)
    dynamic_state_depth_compare_op = int(1000267008)
    dynamic_state_depth_bounds_test_enable = int(1000267009)
    dynamic_state_stencil_test_enable = int(1000267010)
    dynamic_state_stencil_op = int(1000267011)
    dynamic_state_rasterizer_discard_enable = int(1000377001)
    dynamic_state_depth_bias_enable = int(1000377002)
    dynamic_state_primitive_restart_enable = int(1000377004)
    dynamic_state_viewport_w_scaling_nv = int(1000087000)
    dynamic_state_discard_rectangle_ext = int(1000099000)
    dynamic_state_discard_rectangle_enable_ext = int(1000099001)
    dynamic_state_discard_rectangle_mode_ext = int(1000099002)
    dynamic_state_sample_locations_ext = int(1000143000)
    dynamic_state_ray_tracing_pipeline_stack_size_khr = int(1000347000)
    dynamic_state_viewport_shading_rate_palette_nv = int(1000164004)
    dynamic_state_viewport_coarse_sample_order_nv = int(1000164006)
    dynamic_state_exclusive_scissor_enable_nv = int(1000205000)
    dynamic_state_exclusive_scissor_nv = int(1000205001)
    dynamic_state_fragment_shading_rate_khr = int(1000226000)
    dynamic_state_line_stipple_ext = int(1000259000)
    dynamic_state_vertex_input_ext = int(1000352000)
    dynamic_state_patch_control_points_ext = int(1000377000)
    dynamic_state_logic_op_ext = int(1000377003)
    dynamic_state_color_write_enable_ext = int(1000381000)
    dynamic_state_tessellation_domain_origin_ext = int(1000455002)
    dynamic_state_depth_clamp_enable_ext = int(1000455003)
    dynamic_state_polygon_mode_ext = int(1000455004)
    dynamic_state_rasterization_samples_ext = int(1000455005)
    dynamic_state_sample_mask_ext = int(1000455006)
    dynamic_state_alpha_to_coverage_enable_ext = int(1000455007)
    dynamic_state_alpha_to_one_enable_ext = int(1000455008)
    dynamic_state_logic_op_enable_ext = int(1000455009)
    dynamic_state_color_blend_enable_ext = int(1000455010)
    dynamic_state_color_blend_equation_ext = int(1000455011)
    dynamic_state_color_write_mask_ext = int(1000455012)
    dynamic_state_rasterization_stream_ext = int(1000455013)
    dynamic_state_conservative_rasterization_mode_ext = int(1000455014)
    dynamic_state_extra_primitive_overestimation_size_ext = int(1000455015)
    dynamic_state_depth_clip_enable_ext = int(1000455016)
    dynamic_state_sample_locations_enable_ext = int(1000455017)
    dynamic_state_color_blend_advanced_ext = int(1000455018)
    dynamic_state_provoking_vertex_mode_ext = int(1000455019)
    dynamic_state_line_rasterization_mode_ext = int(1000455020)
    dynamic_state_line_stipple_enable_ext = int(1000455021)
    dynamic_state_depth_clip_negative_one_to_one_ext = int(1000455022)
    dynamic_state_viewport_w_scaling_enable_nv = int(1000455023)
    dynamic_state_viewport_swizzle_nv = int(1000455024)
    dynamic_state_coverage_to_color_enable_nv = int(1000455025)
    dynamic_state_coverage_to_color_location_nv = int(1000455026)
    dynamic_state_coverage_modulation_mode_nv = int(1000455027)
    dynamic_state_coverage_modulation_table_enable_nv = int(1000455028)
    dynamic_state_coverage_modulation_table_nv = int(1000455029)
    dynamic_state_shading_rate_image_enable_nv = int(1000455030)
    dynamic_state_representative_fragment_test_enable_nv = int(1000455031)
    dynamic_state_coverage_reduction_mode_nv = int(1000455032)
    dynamic_state_attachment_feedback_loop_enable_ext = int(1000524000)
    dynamic_state_max_enum = int(0x7FFFFFFF)
}


pub enum FrontFace {
    front_face_counter_clockwise = int(0)
    front_face_clockwise = int(1)
    front_face_max_enum = int(0x7FFFFFFF)
}


pub enum VertexInputRate {
    vertex_input_rate_vertex = int(0)
    vertex_input_rate_instance = int(1)
    vertex_input_rate_max_enum = int(0x7FFFFFFF)
}


pub enum PrimitiveTopology {
    primitive_topology_point_list = int(0)
    primitive_topology_line_list = int(1)
    primitive_topology_line_strip = int(2)
    primitive_topology_triangle_list = int(3)
    primitive_topology_triangle_strip = int(4)
    primitive_topology_triangle_fan = int(5)
    primitive_topology_line_list_with_adjacency = int(6)
    primitive_topology_line_strip_with_adjacency = int(7)
    primitive_topology_triangle_list_with_adjacency = int(8)
    primitive_topology_triangle_strip_with_adjacency = int(9)
    primitive_topology_patch_list = int(10)
    primitive_topology_max_enum = int(0x7FFFFFFF)
}


pub enum PolygonMode {
    polygon_mode_fill = int(0)
    polygon_mode_line = int(1)
    polygon_mode_point = int(2)
    polygon_mode_fill_rectangle_nv = int(1000153000)
    polygon_mode_max_enum = int(0x7FFFFFFF)
}


pub enum StencilOp {
    stencil_op_keep = int(0)
    stencil_op_zero = int(1)
    stencil_op_replace = int(2)
    stencil_op_increment_and_clamp = int(3)
    stencil_op_decrement_and_clamp = int(4)
    stencil_op_invert = int(5)
    stencil_op_increment_and_wrap = int(6)
    stencil_op_decrement_and_wrap = int(7)
    stencil_op_max_enum = int(0x7FFFFFFF)
}


pub enum LogicOp {
    logic_op_clear = int(0)
    logic_op_and = int(1)
    logic_op_and_reverse = int(2)
    logic_op_copy = int(3)
    logic_op_and_inverted = int(4)
    logic_op_no_op = int(5)
    logic_op_xor = int(6)
    logic_op_or = int(7)
    logic_op_nor = int(8)
    logic_op_equivalent = int(9)
    logic_op_invert = int(10)
    logic_op_or_reverse = int(11)
    logic_op_copy_inverted = int(12)
    logic_op_or_inverted = int(13)
    logic_op_nand = int(14)
    logic_op_set = int(15)
    logic_op_max_enum = int(0x7FFFFFFF)
}


pub enum BorderColor {
    border_color_float_transparent_black = int(0)
    border_color_int_transparent_black = int(1)
    border_color_float_opaque_black = int(2)
    border_color_int_opaque_black = int(3)
    border_color_float_opaque_white = int(4)
    border_color_int_opaque_white = int(5)
    border_color_float_custom_ext = int(1000287003)
    border_color_int_custom_ext = int(1000287004)
    border_color_max_enum = int(0x7FFFFFFF)
}


pub enum Filter {
    filter_nearest = int(0)
    filter_linear = int(1)
    filter_cubic_ext = int(1000015000)
    filter_max_enum = int(0x7FFFFFFF)
}


pub enum SamplerAddressMode {
    sampler_address_mode_repeat = int(0)
    sampler_address_mode_mirrored_repeat = int(1)
    sampler_address_mode_clamp_to_edge = int(2)
    sampler_address_mode_clamp_to_border = int(3)
    sampler_address_mode_mirror_clamp_to_edge = int(4)
    sampler_address_mode_max_enum = int(0x7FFFFFFF)
}


pub enum SamplerMipmapMode {
    sampler_mipmap_mode_nearest = int(0)
    sampler_mipmap_mode_linear = int(1)
    sampler_mipmap_mode_max_enum = int(0x7FFFFFFF)
}


pub enum DescriptorType {
    descriptor_type_sampler = int(0)
    descriptor_type_combined_image_sampler = int(1)
    descriptor_type_sampled_image = int(2)
    descriptor_type_storage_image = int(3)
    descriptor_type_uniform_texel_buffer = int(4)
    descriptor_type_storage_texel_buffer = int(5)
    descriptor_type_uniform_buffer = int(6)
    descriptor_type_storage_buffer = int(7)
    descriptor_type_uniform_buffer_dynamic = int(8)
    descriptor_type_storage_buffer_dynamic = int(9)
    descriptor_type_input_attachment = int(10)
    descriptor_type_inline_uniform_block = int(1000138000)
    descriptor_type_acceleration_structure_khr = int(1000150000)
    descriptor_type_acceleration_structure_nv = int(1000165000)
    descriptor_type_sample_weight_image_qcom = int(1000440000)
    descriptor_type_block_match_image_qcom = int(1000440001)
    descriptor_type_mutable_ext = int(1000351000)
    descriptor_type_max_enum = int(0x7FFFFFFF)
}


pub enum AttachmentLoadOp {
    attachment_load_op_load = int(0)
    attachment_load_op_clear = int(1)
    attachment_load_op_dont_care = int(2)
    attachment_load_op_none_ext = int(1000400000)
    attachment_load_op_max_enum = int(0x7FFFFFFF)
}


pub enum AttachmentStoreOp {
    attachment_store_op_store = int(0)
    attachment_store_op_dont_care = int(1)
    attachment_store_op_none = int(1000301000)
    attachment_store_op_max_enum = int(0x7FFFFFFF)
}


pub enum PipelineBindPoint {
    pipeline_bind_point_graphics = int(0)
    pipeline_bind_point_compute = int(1)
    pipeline_bind_point_ray_tracing_khr = int(1000165000)
    pipeline_bind_point_subpass_shading_huawei = int(1000369003)
    pipeline_bind_point_max_enum = int(0x7FFFFFFF)
}


pub enum CommandBufferLevel {
    command_buffer_level_primary = int(0)
    command_buffer_level_secondary = int(1)
    command_buffer_level_max_enum = int(0x7FFFFFFF)
}


pub enum IndexType {
    index_type_uint16 = int(0)
    index_type_uint32 = int(1)
    index_type_none_khr = int(1000165000)
    index_type_uint8_ext = int(1000265000)
    index_type_max_enum = int(0x7FFFFFFF)
}


pub enum SubpassContents {
    subpass_contents_inline = int(0)
    subpass_contents_secondary_command_buffers = int(1)
    subpass_contents_inline_and_secondary_command_buffers_ext = int(1000451000)
    subpass_contents_max_enum = int(0x7FFFFFFF)
}


pub enum AccessFlagBits {
    access_indirect_command_read_bit = int(0x00000001)
    access_index_read_bit = int(0x00000002)
    access_vertex_attribute_read_bit = int(0x00000004)
    access_uniform_read_bit = int(0x00000008)
    access_input_attachment_read_bit = int(0x00000010)
    access_shader_read_bit = int(0x00000020)
    access_shader_write_bit = int(0x00000040)
    access_color_attachment_read_bit = int(0x00000080)
    access_color_attachment_write_bit = int(0x00000100)
    access_depth_stencil_attachment_read_bit = int(0x00000200)
    access_depth_stencil_attachment_write_bit = int(0x00000400)
    access_transfer_read_bit = int(0x00000800)
    access_transfer_write_bit = int(0x00001000)
    access_host_read_bit = int(0x00002000)
    access_host_write_bit = int(0x00004000)
    access_memory_read_bit = int(0x00008000)
    access_memory_write_bit = int(0x00010000)
    access_none = int(0)
    access_transform_feedback_write_bit_ext = int(0x02000000)
    access_transform_feedback_counter_read_bit_ext = int(0x04000000)
    access_transform_feedback_counter_write_bit_ext = int(0x08000000)
    access_conditional_rendering_read_bit_ext = int(0x00100000)
    access_color_attachment_read_noncoherent_bit_ext = int(0x00080000)
    access_acceleration_structure_read_bit_khr = int(0x00200000)
    access_acceleration_structure_write_bit_khr = int(0x00400000)
    access_fragment_density_map_read_bit_ext = int(0x01000000)
    access_fragment_shading_rate_attachment_read_bit_khr = int(0x00800000)
    access_command_preprocess_read_bit_nv = int(0x00020000)
    access_command_preprocess_write_bit_nv = int(0x00040000)
    access_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type AccessFlags = u32

pub enum ImageAspectFlagBits {
    image_aspect_color_bit = int(0x00000001)
    image_aspect_depth_bit = int(0x00000002)
    image_aspect_stencil_bit = int(0x00000004)
    image_aspect_metadata_bit = int(0x00000008)
    image_aspect_plane_0_bit = int(0x00000010)
    image_aspect_plane_1_bit = int(0x00000020)
    image_aspect_plane_2_bit = int(0x00000040)
    image_aspect_none = int(0)
    image_aspect_memory_plane_0_bit_ext = int(0x00000080)
    image_aspect_memory_plane_1_bit_ext = int(0x00000100)
    image_aspect_memory_plane_2_bit_ext = int(0x00000200)
    image_aspect_memory_plane_3_bit_ext = int(0x00000400)
    image_aspect_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ImageAspectFlags = u32

pub enum FormatFeatureFlagBits {
    format_feature_sampled_image_bit = int(0x00000001)
    format_feature_storage_image_bit = int(0x00000002)
    format_feature_storage_image_atomic_bit = int(0x00000004)
    format_feature_uniform_texel_buffer_bit = int(0x00000008)
    format_feature_storage_texel_buffer_bit = int(0x00000010)
    format_feature_storage_texel_buffer_atomic_bit = int(0x00000020)
    format_feature_vertex_buffer_bit = int(0x00000040)
    format_feature_color_attachment_bit = int(0x00000080)
    format_feature_color_attachment_blend_bit = int(0x00000100)
    format_feature_depth_stencil_attachment_bit = int(0x00000200)
    format_feature_blit_src_bit = int(0x00000400)
    format_feature_blit_dst_bit = int(0x00000800)
    format_feature_sampled_image_filter_linear_bit = int(0x00001000)
    format_feature_transfer_src_bit = int(0x00004000)
    format_feature_transfer_dst_bit = int(0x00008000)
    format_feature_midpoint_chroma_samples_bit = int(0x00020000)
    format_feature_sampled_image_ycbcr_conversion_linear_filter_bit = int(0x00040000)
    format_feature_sampled_image_ycbcr_conversion_separate_reconstruction_filter_bit = int(0x00080000)
    format_feature_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_bit = int(0x00100000)
    format_feature_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_forceable_bit = int(0x00200000)
    format_feature_disjoint_bit = int(0x00400000)
    format_feature_cosited_chroma_samples_bit = int(0x00800000)
    format_feature_sampled_image_filter_minmax_bit = int(0x00010000)
    format_feature_video_decode_output_bit_khr = int(0x02000000)
    format_feature_video_decode_dpb_bit_khr = int(0x04000000)
    format_feature_acceleration_structure_vertex_buffer_bit_khr = int(0x20000000)
    format_feature_sampled_image_filter_cubic_bit_ext = int(0x00002000)
    format_feature_fragment_density_map_bit_ext = int(0x01000000)
    format_feature_fragment_shading_rate_attachment_bit_khr = int(0x40000000)
    format_feature_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type FormatFeatureFlags = u32

pub enum ImageCreateFlagBits {
    image_create_sparse_binding_bit = int(0x00000001)
    image_create_sparse_residency_bit = int(0x00000002)
    image_create_sparse_aliased_bit = int(0x00000004)
    image_create_mutable_format_bit = int(0x00000008)
    image_create_cube_compatible_bit = int(0x00000010)
    image_create_alias_bit = int(0x00000400)
    image_create_split_instance_bind_regions_bit = int(0x00000040)
    image_create_2d_array_compatible_bit = int(0x00000020)
    image_create_block_texel_view_compatible_bit = int(0x00000080)
    image_create_extended_usage_bit = int(0x00000100)
    image_create_protected_bit = int(0x00000800)
    image_create_disjoint_bit = int(0x00000200)
    image_create_corner_sampled_bit_nv = int(0x00002000)
    image_create_sample_locations_compatible_depth_bit_ext = int(0x00001000)
    image_create_subsampled_bit_ext = int(0x00004000)
    image_create_descriptor_buffer_capture_replay_bit_ext = int(0x00010000)
    image_create_multisampled_render_to_single_sampled_bit_ext = int(0x00040000)
    image_create_2d_view_compatible_bit_ext = int(0x00020000)
    image_create_fragment_density_map_offset_bit_qcom = int(0x00008000)
    image_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ImageCreateFlags = u32

pub enum SampleCountFlagBits {
    sample_count_1_bit = int(0x00000001)
    sample_count_2_bit = int(0x00000002)
    sample_count_4_bit = int(0x00000004)
    sample_count_8_bit = int(0x00000008)
    sample_count_16_bit = int(0x00000010)
    sample_count_32_bit = int(0x00000020)
    sample_count_64_bit = int(0x00000040)
    sample_count_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type SampleCountFlags = u32

pub enum ImageUsageFlagBits {
    image_usage_transfer_src_bit = int(0x00000001)
    image_usage_transfer_dst_bit = int(0x00000002)
    image_usage_sampled_bit = int(0x00000004)
    image_usage_storage_bit = int(0x00000008)
    image_usage_color_attachment_bit = int(0x00000010)
    image_usage_depth_stencil_attachment_bit = int(0x00000020)
    image_usage_transient_attachment_bit = int(0x00000040)
    image_usage_input_attachment_bit = int(0x00000080)
    image_usage_video_decode_dst_bit_khr = int(0x00000400)
    image_usage_video_decode_src_bit_khr = int(0x00000800)
    image_usage_video_decode_dpb_bit_khr = int(0x00001000)
    image_usage_fragment_density_map_bit_ext = int(0x00000200)
    image_usage_fragment_shading_rate_attachment_bit_khr = int(0x00000100)
    image_usage_host_transfer_bit_ext = int(0x00400000)
    image_usage_attachment_feedback_loop_bit_ext = int(0x00080000)
    image_usage_invocation_mask_bit_huawei = int(0x00040000)
    image_usage_sample_weight_bit_qcom = int(0x00100000)
    image_usage_sample_block_match_bit_qcom = int(0x00200000)
    image_usage_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ImageUsageFlags = u32

pub enum InstanceCreateFlagBits {
    instance_create_enumerate_portability_bit_khr = int(0x00000001)
    instance_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type InstanceCreateFlags = u32

pub enum MemoryHeapFlagBits {
    memory_heap_device_local_bit = int(0x00000001)
    memory_heap_multi_instance_bit = int(0x00000002)
    memory_heap_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type MemoryHeapFlags = u32

pub enum MemoryPropertyFlagBits {
    memory_property_device_local_bit = int(0x00000001)
    memory_property_host_visible_bit = int(0x00000002)
    memory_property_host_coherent_bit = int(0x00000004)
    memory_property_host_cached_bit = int(0x00000008)
    memory_property_lazily_allocated_bit = int(0x00000010)
    memory_property_protected_bit = int(0x00000020)
    memory_property_device_coherent_bit_amd = int(0x00000040)
    memory_property_device_uncached_bit_amd = int(0x00000080)
    memory_property_rdma_capable_bit_nv = int(0x00000100)
    memory_property_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type MemoryPropertyFlags = u32

pub enum QueueFlagBits {
    queue_graphics_bit = int(0x00000001)
    queue_compute_bit = int(0x00000002)
    queue_transfer_bit = int(0x00000004)
    queue_sparse_binding_bit = int(0x00000008)
    queue_protected_bit = int(0x00000010)
    queue_video_decode_bit_khr = int(0x00000020)
    queue_optical_flow_bit_nv = int(0x00000100)
    queue_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type QueueFlags = u32
pub type DeviceCreateFlags = u32

pub enum DeviceQueueCreateFlagBits {
    device_queue_create_protected_bit = int(0x00000001)
    device_queue_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type DeviceQueueCreateFlags = u32

pub enum PipelineStageFlagBits {
    pipeline_stage_top_of_pipe_bit = int(0x00000001)
    pipeline_stage_draw_indirect_bit = int(0x00000002)
    pipeline_stage_vertex_input_bit = int(0x00000004)
    pipeline_stage_vertex_shader_bit = int(0x00000008)
    pipeline_stage_tessellation_control_shader_bit = int(0x00000010)
    pipeline_stage_tessellation_evaluation_shader_bit = int(0x00000020)
    pipeline_stage_geometry_shader_bit = int(0x00000040)
    pipeline_stage_fragment_shader_bit = int(0x00000080)
    pipeline_stage_early_fragment_tests_bit = int(0x00000100)
    pipeline_stage_late_fragment_tests_bit = int(0x00000200)
    pipeline_stage_color_attachment_output_bit = int(0x00000400)
    pipeline_stage_compute_shader_bit = int(0x00000800)
    pipeline_stage_transfer_bit = int(0x00001000)
    pipeline_stage_bottom_of_pipe_bit = int(0x00002000)
    pipeline_stage_host_bit = int(0x00004000)
    pipeline_stage_all_graphics_bit = int(0x00008000)
    pipeline_stage_all_commands_bit = int(0x00010000)
    pipeline_stage_none = int(0)
    pipeline_stage_transform_feedback_bit_ext = int(0x01000000)
    pipeline_stage_conditional_rendering_bit_ext = int(0x00040000)
    pipeline_stage_acceleration_structure_build_bit_khr = int(0x02000000)
    pipeline_stage_ray_tracing_shader_bit_khr = int(0x00200000)
    pipeline_stage_fragment_density_process_bit_ext = int(0x00800000)
    pipeline_stage_fragment_shading_rate_attachment_bit_khr = int(0x00400000)
    pipeline_stage_command_preprocess_bit_nv = int(0x00020000)
    pipeline_stage_task_shader_bit_ext = int(0x00080000)
    pipeline_stage_mesh_shader_bit_ext = int(0x00100000)
    pipeline_stage_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type PipelineStageFlags = u32
pub type MemoryMapFlags = u32

pub enum SparseMemoryBindFlagBits {
    sparse_memory_bind_metadata_bit = int(0x00000001)
    sparse_memory_bind_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type SparseMemoryBindFlags = u32

pub enum SparseImageFormatFlagBits {
    sparse_image_format_single_miptail_bit = int(0x00000001)
    sparse_image_format_aligned_mip_size_bit = int(0x00000002)
    sparse_image_format_nonstandard_block_size_bit = int(0x00000004)
    sparse_image_format_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type SparseImageFormatFlags = u32

pub enum FenceCreateFlagBits {
    fence_create_signaled_bit = int(0x00000001)
    fence_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type FenceCreateFlags = u32
pub type SemaphoreCreateFlags = u32

pub enum EventCreateFlagBits {
    event_create_device_only_bit = int(0x00000001)
    event_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type EventCreateFlags = u32

pub enum QueryPipelineStatisticFlagBits {
    query_pipeline_statistic_input_assembly_vertices_bit = int(0x00000001)
    query_pipeline_statistic_input_assembly_primitives_bit = int(0x00000002)
    query_pipeline_statistic_vertex_shader_invocations_bit = int(0x00000004)
    query_pipeline_statistic_geometry_shader_invocations_bit = int(0x00000008)
    query_pipeline_statistic_geometry_shader_primitives_bit = int(0x00000010)
    query_pipeline_statistic_clipping_invocations_bit = int(0x00000020)
    query_pipeline_statistic_clipping_primitives_bit = int(0x00000040)
    query_pipeline_statistic_fragment_shader_invocations_bit = int(0x00000080)
    query_pipeline_statistic_tessellation_control_shader_patches_bit = int(0x00000100)
    query_pipeline_statistic_tessellation_evaluation_shader_invocations_bit = int(0x00000200)
    query_pipeline_statistic_compute_shader_invocations_bit = int(0x00000400)
    query_pipeline_statistic_task_shader_invocations_bit_ext = int(0x00000800)
    query_pipeline_statistic_mesh_shader_invocations_bit_ext = int(0x00001000)
    query_pipeline_statistic_cluster_culling_shader_invocations_bit_huawei = int(0x00002000)
    query_pipeline_statistic_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type QueryPipelineStatisticFlags = u32
pub type QueryPoolCreateFlags = u32

pub enum QueryResultFlagBits {
    query_result_64_bit = int(0x00000001)
    query_result_wait_bit = int(0x00000002)
    query_result_with_availability_bit = int(0x00000004)
    query_result_partial_bit = int(0x00000008)
    query_result_with_status_bit_khr = int(0x00000010)
    query_result_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type QueryResultFlags = u32

pub enum BufferCreateFlagBits {
    buffer_create_sparse_binding_bit = int(0x00000001)
    buffer_create_sparse_residency_bit = int(0x00000002)
    buffer_create_sparse_aliased_bit = int(0x00000004)
    buffer_create_protected_bit = int(0x00000008)
    buffer_create_device_address_capture_replay_bit = int(0x00000010)
    buffer_create_descriptor_buffer_capture_replay_bit_ext = int(0x00000020)
    buffer_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type BufferCreateFlags = u32

pub enum BufferUsageFlagBits {
    buffer_usage_transfer_src_bit = int(0x00000001)
    buffer_usage_transfer_dst_bit = int(0x00000002)
    buffer_usage_uniform_texel_buffer_bit = int(0x00000004)
    buffer_usage_storage_texel_buffer_bit = int(0x00000008)
    buffer_usage_uniform_buffer_bit = int(0x00000010)
    buffer_usage_storage_buffer_bit = int(0x00000020)
    buffer_usage_index_buffer_bit = int(0x00000040)
    buffer_usage_vertex_buffer_bit = int(0x00000080)
    buffer_usage_indirect_buffer_bit = int(0x00000100)
    buffer_usage_shader_device_address_bit = int(0x00020000)
    buffer_usage_video_decode_src_bit_khr = int(0x00002000)
    buffer_usage_video_decode_dst_bit_khr = int(0x00004000)
    buffer_usage_transform_feedback_buffer_bit_ext = int(0x00000800)
    buffer_usage_transform_feedback_counter_buffer_bit_ext = int(0x00001000)
    buffer_usage_conditional_rendering_bit_ext = int(0x00000200)
    buffer_usage_acceleration_structure_build_input_read_only_bit_khr = int(0x00080000)
    buffer_usage_acceleration_structure_storage_bit_khr = int(0x00100000)
    buffer_usage_shader_binding_table_bit_khr = int(0x00000400)
    buffer_usage_sampler_descriptor_buffer_bit_ext = int(0x00200000)
    buffer_usage_resource_descriptor_buffer_bit_ext = int(0x00400000)
    buffer_usage_push_descriptors_descriptor_buffer_bit_ext = int(0x04000000)
    buffer_usage_micromap_build_input_read_only_bit_ext = int(0x00800000)
    buffer_usage_micromap_storage_bit_ext = int(0x01000000)
    buffer_usage_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type BufferUsageFlags = u32
pub type BufferViewCreateFlags = u32

pub enum ImageViewCreateFlagBits {
    image_view_create_fragment_density_map_dynamic_bit_ext = int(0x00000001)
    image_view_create_descriptor_buffer_capture_replay_bit_ext = int(0x00000004)
    image_view_create_fragment_density_map_deferred_bit_ext = int(0x00000002)
    image_view_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ImageViewCreateFlags = u32
pub type ShaderModuleCreateFlags = u32

pub enum PipelineCacheCreateFlagBits {
    pipeline_cache_create_externally_synchronized_bit = int(0x00000001)
    pipeline_cache_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type PipelineCacheCreateFlags = u32

pub enum ColorComponentFlagBits {
    color_component_r_bit = int(0x00000001)
    color_component_g_bit = int(0x00000002)
    color_component_b_bit = int(0x00000004)
    color_component_a_bit = int(0x00000008)
    color_component_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ColorComponentFlags = u32

pub enum PipelineCreateFlagBits {
    pipeline_create_disable_optimization_bit = int(0x00000001)
    pipeline_create_allow_derivatives_bit = int(0x00000002)
    pipeline_create_derivative_bit = int(0x00000004)
    pipeline_create_view_index_from_device_index_bit = int(0x00000008)
    pipeline_create_dispatch_base_bit = int(0x00000010)
    pipeline_create_fail_on_pipeline_compile_required_bit = int(0x00000100)
    pipeline_create_early_return_on_failure_bit = int(0x00000200)
    pipeline_create_rendering_fragment_shading_rate_attachment_bit_khr = int(0x00200000)
    pipeline_create_rendering_fragment_density_map_attachment_bit_ext = int(0x00400000)
    pipeline_create_ray_tracing_no_null_any_hit_shaders_bit_khr = int(0x00004000)
    pipeline_create_ray_tracing_no_null_closest_hit_shaders_bit_khr = int(0x00008000)
    pipeline_create_ray_tracing_no_null_miss_shaders_bit_khr = int(0x00010000)
    pipeline_create_ray_tracing_no_null_intersection_shaders_bit_khr = int(0x00020000)
    pipeline_create_ray_tracing_skip_triangles_bit_khr = int(0x00001000)
    pipeline_create_ray_tracing_skip_aabbs_bit_khr = int(0x00002000)
    pipeline_create_ray_tracing_shader_group_handle_capture_replay_bit_khr = int(0x00080000)
    pipeline_create_defer_compile_bit_nv = int(0x00000020)
    pipeline_create_capture_statistics_bit_khr = int(0x00000040)
    pipeline_create_capture_internal_representations_bit_khr = int(0x00000080)
    pipeline_create_indirect_bindable_bit_nv = int(0x00040000)
    pipeline_create_library_bit_khr = int(0x00000800)
    pipeline_create_descriptor_buffer_bit_ext = int(0x20000000)
    pipeline_create_retain_link_time_optimization_info_bit_ext = int(0x00800000)
    pipeline_create_link_time_optimization_bit_ext = int(0x00000400)
    pipeline_create_ray_tracing_allow_motion_bit_nv = int(0x00100000)
    pipeline_create_color_attachment_feedback_loop_bit_ext = int(0x02000000)
    pipeline_create_depth_stencil_attachment_feedback_loop_bit_ext = int(0x04000000)
    pipeline_create_ray_tracing_opacity_micromap_bit_ext = int(0x01000000)
    pipeline_create_no_protected_access_bit_ext = int(0x08000000)
    pipeline_create_protected_access_only_bit_ext = int(0x40000000)
    pipeline_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type PipelineCreateFlags = u32

pub enum PipelineShaderStageCreateFlagBits {
    pipeline_shader_stage_create_allow_varying_subgroup_size_bit = int(0x00000001)
    pipeline_shader_stage_create_require_full_subgroups_bit = int(0x00000002)
    pipeline_shader_stage_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type PipelineShaderStageCreateFlags = u32

pub enum ShaderStageFlagBits {
    shader_stage_vertex_bit = int(0x00000001)
    shader_stage_tessellation_control_bit = int(0x00000002)
    shader_stage_tessellation_evaluation_bit = int(0x00000004)
    shader_stage_geometry_bit = int(0x00000008)
    shader_stage_fragment_bit = int(0x00000010)
    shader_stage_compute_bit = int(0x00000020)
    shader_stage_all_graphics = int(0x0000001F)
    shader_stage_all = int(0x7FFFFFFF)
    shader_stage_raygen_bit_khr = int(0x00000100)
    shader_stage_any_hit_bit_khr = int(0x00000200)
    shader_stage_closest_hit_bit_khr = int(0x00000400)
    shader_stage_miss_bit_khr = int(0x00000800)
    shader_stage_intersection_bit_khr = int(0x00001000)
    shader_stage_callable_bit_khr = int(0x00002000)
    shader_stage_task_bit_ext = int(0x00000040)
    shader_stage_mesh_bit_ext = int(0x00000080)
    shader_stage_subpass_shading_bit_huawei = int(0x00004000)
    shader_stage_cluster_culling_bit_huawei = int(0x00080000)
    shader_stage_flag_bits_max_enum = int(0x7FFFFFFF)
}


pub enum CullModeFlagBits {
    cull_mode_none = int(0)
    cull_mode_front_bit = int(0x00000001)
    cull_mode_back_bit = int(0x00000002)
    cull_mode_front_and_back = int(0x00000003)
    cull_mode_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type CullModeFlags = u32
pub type PipelineVertexInputStateCreateFlags = u32
pub type PipelineInputAssemblyStateCreateFlags = u32
pub type PipelineTessellationStateCreateFlags = u32
pub type PipelineViewportStateCreateFlags = u32
pub type PipelineRasterizationStateCreateFlags = u32
pub type PipelineMultisampleStateCreateFlags = u32

pub enum PipelineDepthStencilStateCreateFlagBits {
    pipeline_depth_stencil_state_create_rasterization_order_attachment_depth_access_bit_ext = int(0x00000001)
    pipeline_depth_stencil_state_create_rasterization_order_attachment_stencil_access_bit_ext = int(0x00000002)
    pipeline_depth_stencil_state_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type PipelineDepthStencilStateCreateFlags = u32

pub enum PipelineColorBlendStateCreateFlagBits {
    pipeline_color_blend_state_create_rasterization_order_attachment_access_bit_ext = int(0x00000001)
    pipeline_color_blend_state_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type PipelineColorBlendStateCreateFlags = u32
pub type PipelineDynamicStateCreateFlags = u32

pub enum PipelineLayoutCreateFlagBits {
    pipeline_layout_create_independent_sets_bit_ext = int(0x00000002)
    pipeline_layout_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type PipelineLayoutCreateFlags = u32
pub type ShaderStageFlags = u32

pub enum SamplerCreateFlagBits {
    sampler_create_subsampled_bit_ext = int(0x00000001)
    sampler_create_subsampled_coarse_reconstruction_bit_ext = int(0x00000002)
    sampler_create_descriptor_buffer_capture_replay_bit_ext = int(0x00000008)
    sampler_create_non_seamless_cube_map_bit_ext = int(0x00000004)
    sampler_create_image_processing_bit_qcom = int(0x00000010)
    sampler_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type SamplerCreateFlags = u32

pub enum DescriptorPoolCreateFlagBits {
    descriptor_pool_create_free_descriptor_set_bit = int(0x00000001)
    descriptor_pool_create_update_after_bind_bit = int(0x00000002)
    descriptor_pool_create_host_only_bit_ext = int(0x00000004)
    descriptor_pool_create_allow_overallocation_sets_bit_nv = int(0x00000008)
    descriptor_pool_create_allow_overallocation_pools_bit_nv = int(0x00000010)
    descriptor_pool_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type DescriptorPoolCreateFlags = u32
pub type DescriptorPoolResetFlags = u32

pub enum DescriptorSetLayoutCreateFlagBits {
    descriptor_set_layout_create_update_after_bind_pool_bit = int(0x00000002)
    descriptor_set_layout_create_push_descriptor_bit_khr = int(0x00000001)
    descriptor_set_layout_create_descriptor_buffer_bit_ext = int(0x00000010)
    descriptor_set_layout_create_embedded_immutable_samplers_bit_ext = int(0x00000020)
    descriptor_set_layout_create_indirect_bindable_bit_nv = int(0x00000080)
    descriptor_set_layout_create_host_only_pool_bit_ext = int(0x00000004)
    descriptor_set_layout_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type DescriptorSetLayoutCreateFlags = u32

pub enum AttachmentDescriptionFlagBits {
    attachment_description_may_alias_bit = int(0x00000001)
    attachment_description_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type AttachmentDescriptionFlags = u32

pub enum DependencyFlagBits {
    dependency_by_region_bit = int(0x00000001)
    dependency_device_group_bit = int(0x00000004)
    dependency_view_local_bit = int(0x00000002)
    dependency_feedback_loop_bit_ext = int(0x00000008)
    dependency_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type DependencyFlags = u32

pub enum FramebufferCreateFlagBits {
    framebuffer_create_imageless_bit = int(0x00000001)
    framebuffer_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type FramebufferCreateFlags = u32

pub enum RenderPassCreateFlagBits {
    render_pass_create_transform_bit_qcom = int(0x00000002)
    render_pass_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type RenderPassCreateFlags = u32

pub enum SubpassDescriptionFlagBits {
    subpass_description_per_view_attributes_bit_nvx = int(0x00000001)
    subpass_description_per_view_position_x_only_bit_nvx = int(0x00000002)
    subpass_description_fragment_region_bit_qcom = int(0x00000004)
    subpass_description_shader_resolve_bit_qcom = int(0x00000008)
    subpass_description_rasterization_order_attachment_color_access_bit_ext = int(0x00000010)
    subpass_description_rasterization_order_attachment_depth_access_bit_ext = int(0x00000020)
    subpass_description_rasterization_order_attachment_stencil_access_bit_ext = int(0x00000040)
    subpass_description_enable_legacy_dithering_bit_ext = int(0x00000080)
    subpass_description_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type SubpassDescriptionFlags = u32

pub enum CommandPoolCreateFlagBits {
    command_pool_create_transient_bit = int(0x00000001)
    command_pool_create_reset_command_buffer_bit = int(0x00000002)
    command_pool_create_protected_bit = int(0x00000004)
    command_pool_create_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type CommandPoolCreateFlags = u32

pub enum CommandPoolResetFlagBits {
    command_pool_reset_release_resources_bit = int(0x00000001)
    command_pool_reset_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type CommandPoolResetFlags = u32

pub enum CommandBufferUsageFlagBits {
    command_buffer_usage_one_time_submit_bit = int(0x00000001)
    command_buffer_usage_render_pass_continue_bit = int(0x00000002)
    command_buffer_usage_simultaneous_use_bit = int(0x00000004)
    command_buffer_usage_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type CommandBufferUsageFlags = u32

pub enum QueryControlFlagBits {
    query_control_precise_bit = int(0x00000001)
    query_control_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type QueryControlFlags = u32

pub enum CommandBufferResetFlagBits {
    command_buffer_reset_release_resources_bit = int(0x00000001)
    command_buffer_reset_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type CommandBufferResetFlags = u32

pub enum StencilFaceFlagBits {
    stencil_face_front_bit = int(0x00000001)
    stencil_face_back_bit = int(0x00000002)
    stencil_face_front_and_back = int(0x00000003)
    stencil_face_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type StencilFaceFlags = u32
pub struct Extent2D {
mut:
    width           u32
    height          u32
} 

pub struct Extent3D {
mut:
    width           u32
    height          u32
    depth           u32
} 

pub struct Offset2D {
mut:
    x              i32
    y              i32
} 

pub struct Offset3D {
mut:
    x              i32
    y              i32
    z              i32
} 

pub struct Rect2D {
mut:
    offset            Offset2D
    extent            Extent2D
} 

pub struct BaseInStructure {
mut:
    s_type                                 StructureType
    p_next                                 &BaseInStructure
} 

pub struct BaseOutStructure {
mut:
    s_type                            StructureType
    p_next                            &BaseOutStructure
} 

pub struct BufferMemoryBarrier {
mut:
    s_type                 StructureType
    p_next                 voidptr
    src_access_mask        AccessFlags
    dst_access_mask        AccessFlags
    src_queue_family_index u32
    dst_queue_family_index u32
    buffer                 C.Buffer
    offset                 DeviceSize
    size                   DeviceSize
} 

pub struct DispatchIndirectCommand {
mut:
    x               u32
    y               u32
    z               u32
} 

pub struct DrawIndexedIndirectCommand {
mut:
    index_count     u32
    instance_count  u32
    first_index     u32
    vertex_offset   i32
    first_instance  u32
} 

pub struct DrawIndirectCommand {
mut:
    vertex_count    u32
    instance_count  u32
    first_vertex    u32
    first_instance  u32
} 

pub struct ImageSubresourceRange {
mut:
    aspect_mask               ImageAspectFlags
    base_mip_level            u32
    level_count               u32
    base_array_layer          u32
    layer_count               u32
} 

pub struct ImageMemoryBarrier {
mut:
    s_type                         StructureType
    p_next                         voidptr
    src_access_mask                AccessFlags
    dst_access_mask                AccessFlags
    old_layout                     ImageLayout
    new_layout                     ImageLayout
    src_queue_family_index         u32
    dst_queue_family_index         u32
    image                          C.Image
    subresource_range              ImageSubresourceRange
} 

pub struct MemoryBarrier {
mut:
    s_type                 StructureType
    p_next                 voidptr
    src_access_mask        AccessFlags
    dst_access_mask        AccessFlags
} 

pub struct PipelineCacheHeaderVersionOne {
mut:
    header_size                         u32
    header_version                      PipelineCacheHeaderVersion
    vendor_id                           u32
    device_id                           u32
    pipeline_cache_uuid                 []u8
} 

pub type PFN_vkAllocationFunction = fn (   pUserData                         voidptr,   size                              usize,   alignment                         usize,   allocationScope                   SystemAllocationScope) voidptr
pub type PFN_vkFreeFunction = fn (   pUserData                         voidptr,   pMemory                           voidptr) voidptr
pub type PFN_vkInternalAllocationNotification = fn (   pUserData                         voidptr,   size                              usize,   allocationType                    InternalAllocationType,   allocationScope                   SystemAllocationScope) voidptr
pub type PFN_vkInternalFreeNotification = fn (   pUserData                         voidptr,   size                              usize,   allocationType                    InternalAllocationType,   allocationScope                   SystemAllocationScope) voidptr
pub type PFN_vkReallocationFunction = fn (   pUserData                         voidptr,   pOriginal                         voidptr,   size                              usize,   alignment                         usize,   allocationScope                   SystemAllocationScope) voidptr
pub type PFN_vkVoidFunction = fn () 
pub struct AllocationCallbacks {
mut:
    p_user_data                                 voidptr
    pfn_allocation                              PFN_vkAllocationFunction = unsafe { nil }
    pfn_reallocation                            PFN_vkReallocationFunction = unsafe { nil }
    pfn_free                                    PFN_vkFreeFunction = unsafe { nil }
    pfn_internal_allocation                     PFN_vkInternalAllocationNotification = unsafe { nil }
    pfn_internal_free                           PFN_vkInternalFreeNotification = unsafe { nil }
} 

pub struct ApplicationInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    p_application_name     &char
    application_version    u32
    p_engine_name          &char
    engine_version         u32
    api_version            u32
} 

pub struct FormatProperties {
mut:
    linear_tiling_features      FormatFeatureFlags
    optimal_tiling_features     FormatFeatureFlags
    buffer_features             FormatFeatureFlags
} 

pub struct ImageFormatProperties {
mut:
    max_extent                Extent3D
    max_mip_levels            u32
    max_array_layers          u32
    sample_counts             SampleCountFlags
    max_resource_size         DeviceSize
} 

pub struct InstanceCreateInfo {
mut:
    s_type                          StructureType
    p_next                          voidptr
    flags                           InstanceCreateFlags
    p_application_info              &ApplicationInfo
    enabled_layer_count             u32
    pp_enabled_layer_names          &char
    enabled_extension_count         u32
    pp_enabled_extension_names      &char
} 

pub struct MemoryHeap {
mut:
    size                     DeviceSize
    flags                    MemoryHeapFlags
} 

pub struct MemoryType {
mut:
    property_flags               MemoryPropertyFlags
    heap_index                   u32
} 

pub struct PhysicalDeviceFeatures {
mut:
    robust_buffer_access Bool32
    full_draw_index_uint32 Bool32
    image_cube_array Bool32
    independent_blend Bool32
    geometry_shader Bool32
    tessellation_shader Bool32
    sample_rate_shading Bool32
    dual_src_blend  Bool32
    logic_op        Bool32
    multi_draw_indirect Bool32
    draw_indirect_first_instance Bool32
    depth_clamp     Bool32
    depth_bias_clamp Bool32
    fill_mode_non_solid Bool32
    depth_bounds    Bool32
    wide_lines      Bool32
    large_points    Bool32
    alpha_to_one    Bool32
    multi_viewport  Bool32
    sampler_anisotropy Bool32
    texture_compression_etc2 Bool32
    texture_compression_astc_ldr Bool32
    texture_compression_bc Bool32
    occlusion_query_precise Bool32
    pipeline_statistics_query Bool32
    vertex_pipeline_stores_and_atomics Bool32
    fragment_stores_and_atomics Bool32
    shader_tessellation_and_geometry_point_size Bool32
    shader_image_gather_extended Bool32
    shader_storage_image_extended_formats Bool32
    shader_storage_image_multisample Bool32
    shader_storage_image_read_without_format Bool32
    shader_storage_image_write_without_format Bool32
    shader_uniform_buffer_array_dynamic_indexing Bool32
    shader_sampled_image_array_dynamic_indexing Bool32
    shader_storage_buffer_array_dynamic_indexing Bool32
    shader_storage_image_array_dynamic_indexing Bool32
    shader_clip_distance Bool32
    shader_cull_distance Bool32
    shader_float64  Bool32
    shader_int64    Bool32
    shader_int16    Bool32
    shader_resource_residency Bool32
    shader_resource_min_lod Bool32
    sparse_binding  Bool32
    sparse_residency_buffer Bool32
    sparse_residency_image2_d Bool32
    sparse_residency_image3_d Bool32
    sparse_residency2_samples Bool32
    sparse_residency4_samples Bool32
    sparse_residency8_samples Bool32
    sparse_residency16_samples Bool32
    sparse_residency_aliased Bool32
    variable_multisample_rate Bool32
    inherited_queries Bool32
} 

pub struct PhysicalDeviceLimits {
mut:
    max_image_dimension1_d    u32
    max_image_dimension2_d    u32
    max_image_dimension3_d    u32
    max_image_dimension_cube  u32
    max_image_array_layers    u32
    max_texel_buffer_elements u32
    max_uniform_buffer_range  u32
    max_storage_buffer_range  u32
    max_push_constants_size   u32
    max_memory_allocation_count u32
    max_sampler_allocation_count u32
    buffer_image_granularity  DeviceSize
    sparse_address_space_size DeviceSize
    max_bound_descriptor_sets u32
    max_per_stage_descriptor_samplers u32
    max_per_stage_descriptor_uniform_buffers u32
    max_per_stage_descriptor_storage_buffers u32
    max_per_stage_descriptor_sampled_images u32
    max_per_stage_descriptor_storage_images u32
    max_per_stage_descriptor_input_attachments u32
    max_per_stage_resources   u32
    max_descriptor_set_samplers u32
    max_descriptor_set_uniform_buffers u32
    max_descriptor_set_uniform_buffers_dynamic u32
    max_descriptor_set_storage_buffers u32
    max_descriptor_set_storage_buffers_dynamic u32
    max_descriptor_set_sampled_images u32
    max_descriptor_set_storage_images u32
    max_descriptor_set_input_attachments u32
    max_vertex_input_attributes u32
    max_vertex_input_bindings u32
    max_vertex_input_attribute_offset u32
    max_vertex_input_binding_stride u32
    max_vertex_output_components u32
    max_tessellation_generation_level u32
    max_tessellation_patch_size u32
    max_tessellation_control_per_vertex_input_components u32
    max_tessellation_control_per_vertex_output_components u32
    max_tessellation_control_per_patch_output_components u32
    max_tessellation_control_total_output_components u32
    max_tessellation_evaluation_input_components u32
    max_tessellation_evaluation_output_components u32
    max_geometry_shader_invocations u32
    max_geometry_input_components u32
    max_geometry_output_components u32
    max_geometry_output_vertices u32
    max_geometry_total_output_components u32
    max_fragment_input_components u32
    max_fragment_output_attachments u32
    max_fragment_dual_src_attachments u32
    max_fragment_combined_output_resources u32
    max_compute_shared_memory_size u32
    max_compute_work_group_count []u32
    max_compute_work_group_invocations u32
    max_compute_work_group_size []u32
    sub_pixel_precision_bits  u32
    sub_texel_precision_bits  u32
    mipmap_precision_bits     u32
    max_draw_indexed_index_value u32
    max_draw_indirect_count   u32
    max_sampler_lod_bias      f32
    max_sampler_anisotropy    f32
    max_viewports             u32
    max_viewport_dimensions   []u32
    viewport_bounds_range     []f32
    viewport_sub_pixel_bits   u32
    min_memory_map_alignment  usize
    min_texel_buffer_offset_alignment DeviceSize
    min_uniform_buffer_offset_alignment DeviceSize
    min_storage_buffer_offset_alignment DeviceSize
    min_texel_offset          i32
    max_texel_offset          u32
    min_texel_gather_offset   i32
    max_texel_gather_offset   u32
    min_interpolation_offset  f32
    max_interpolation_offset  f32
    sub_pixel_interpolation_offset_bits u32
    max_framebuffer_width     u32
    max_framebuffer_height    u32
    max_framebuffer_layers    u32
    framebuffer_color_sample_counts SampleCountFlags
    framebuffer_depth_sample_counts SampleCountFlags
    framebuffer_stencil_sample_counts SampleCountFlags
    framebuffer_no_attachments_sample_counts SampleCountFlags
    max_color_attachments     u32
    sampled_image_color_sample_counts SampleCountFlags
    sampled_image_integer_sample_counts SampleCountFlags
    sampled_image_depth_sample_counts SampleCountFlags
    sampled_image_stencil_sample_counts SampleCountFlags
    storage_image_sample_counts SampleCountFlags
    max_sample_mask_words     u32
    timestamp_compute_and_graphics Bool32
    timestamp_period          f32
    max_clip_distances        u32
    max_cull_distances        u32
    max_combined_clip_and_cull_distances u32
    discrete_queue_priorities u32
    point_size_range          []f32
    line_width_range          []f32
    point_size_granularity    f32
    line_width_granularity    f32
    strict_lines              Bool32
    standard_sample_locations Bool32
    optimal_buffer_copy_offset_alignment DeviceSize
    optimal_buffer_copy_row_pitch_alignment DeviceSize
    non_coherent_atom_size    DeviceSize
} 

pub struct PhysicalDeviceMemoryProperties {
mut:
    memory_type_count   u32
    memory_types        []MemoryType
    memory_heap_count   u32
    memory_heaps        []MemoryHeap
} 

pub struct PhysicalDeviceSparseProperties {
mut:
    residency_standard2_d_block_shape Bool32
    residency_standard2_d_multisample_block_shape Bool32
    residency_standard3_d_block_shape Bool32
    residency_aligned_mip_size Bool32
    residency_non_resident_strict Bool32
} 

pub struct PhysicalDeviceProperties {
mut:
    api_version                             u32
    driver_version                          u32
    vendor_id                               u32
    device_id                               u32
    device_type                             PhysicalDeviceType
    device_name                             []char
    pipeline_cache_uuid                     []u8
    limits                                  PhysicalDeviceLimits
    sparse_properties                       PhysicalDeviceSparseProperties
} 

pub struct QueueFamilyProperties {
mut:
    queue_flags         QueueFlags
    queue_count         u32
    timestamp_valid_bits u32
    min_image_transfer_granularity Extent3D
} 

pub struct DeviceQueueCreateInfo {
mut:
    s_type                          StructureType
    p_next                          voidptr
    flags                           DeviceQueueCreateFlags
    queue_family_index              u32
    queue_count                     u32
    p_queue_priorities              &f32
} 

pub struct DeviceCreateInfo {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    flags                                  DeviceCreateFlags
    queue_create_info_count                u32
    p_queue_create_infos                   &DeviceQueueCreateInfo
    enabled_layer_count                    u32
    pp_enabled_layer_names                 &char
    enabled_extension_count                u32
    pp_enabled_extension_names             &char
    p_enabled_features                     &PhysicalDeviceFeatures
} 

pub struct ExtensionProperties {
mut:
    extension_name  []char
    spec_version    u32
} 

pub struct LayerProperties {
mut:
    layer_name      []char
    spec_version    u32
    implementation_version u32
    description     []char
} 

pub struct SubmitInfo {
mut:
    s_type                             StructureType
    p_next                             voidptr
    wait_semaphore_count               u32
    p_wait_semaphores                  &C.Semaphore
    p_wait_dst_stage_mask              &PipelineStageFlags
    command_buffer_count               u32
    p_command_buffers                  &C.CommandBuffer
    signal_semaphore_count             u32
    p_signal_semaphores                &C.Semaphore
} 

pub struct MappedMemoryRange {
mut:
    s_type                 StructureType
    p_next                 voidptr
    memory                 C.DeviceMemory
    offset                 DeviceSize
    size                   DeviceSize
} 

pub struct MemoryAllocateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    allocation_size        DeviceSize
    memory_type_index      u32
} 

pub struct MemoryRequirements {
mut:
    size                DeviceSize
    alignment           DeviceSize
    memory_type_bits    u32
} 

pub struct SparseMemoryBind {
mut:
    resource_offset                DeviceSize
    size                           DeviceSize
    memory                         C.DeviceMemory
    memory_offset                  DeviceSize
    flags                          SparseMemoryBindFlags
} 

pub struct SparseBufferMemoryBindInfo {
mut:
    buffer                           C.Buffer
    bind_count                       u32
    p_binds                          &SparseMemoryBind
} 

pub struct SparseImageOpaqueMemoryBindInfo {
mut:
    image                            C.Image
    bind_count                       u32
    p_binds                          &SparseMemoryBind
} 

pub struct ImageSubresource {
mut:
    aspect_mask               ImageAspectFlags
    mip_level                 u32
    array_layer               u32
} 

pub struct SparseImageMemoryBind {
mut:
    subresource                    ImageSubresource
    offset                         Offset3D
    extent                         Extent3D
    memory                         C.DeviceMemory
    memory_offset                  DeviceSize
    flags                          SparseMemoryBindFlags
} 

pub struct SparseImageMemoryBindInfo {
mut:
    image                                 C.Image
    bind_count                            u32
    p_binds                               &SparseImageMemoryBind
} 

pub struct BindSparseInfo {
mut:
    s_type                                          StructureType
    p_next                                          voidptr
    wait_semaphore_count                            u32
    p_wait_semaphores                               &C.Semaphore
    buffer_bind_count                               u32
    p_buffer_binds                                  &SparseBufferMemoryBindInfo
    image_opaque_bind_count                         u32
    p_image_opaque_binds                            &SparseImageOpaqueMemoryBindInfo
    image_bind_count                                u32
    p_image_binds                                   &SparseImageMemoryBindInfo
    signal_semaphore_count                          u32
    p_signal_semaphores                             &C.Semaphore
} 

pub struct SparseImageFormatProperties {
mut:
    aspect_mask                     ImageAspectFlags
    image_granularity               Extent3D
    flags                           SparseImageFormatFlags
} 

pub struct SparseImageMemoryRequirements {
mut:
    format_properties                    SparseImageFormatProperties
    image_mip_tail_first_lod             u32
    image_mip_tail_size                  DeviceSize
    image_mip_tail_offset                DeviceSize
    image_mip_tail_stride                DeviceSize
} 

pub struct FenceCreateInfo {
mut:
    s_type                    StructureType
    p_next                    voidptr
    flags                     FenceCreateFlags
} 

pub struct SemaphoreCreateInfo {
mut:
    s_type                        StructureType
    p_next                        voidptr
    flags                         SemaphoreCreateFlags
} 

pub struct EventCreateInfo {
mut:
    s_type                    StructureType
    p_next                    voidptr
    flags                     EventCreateFlags
} 

pub struct QueryPoolCreateInfo {
mut:
    s_type                               StructureType
    p_next                               voidptr
    flags                                QueryPoolCreateFlags
    query_type                           QueryType
    query_count                          u32
    pipeline_statistics                  QueryPipelineStatisticFlags
} 

pub struct BufferCreateInfo {
mut:
    s_type                     StructureType
    p_next                     voidptr
    flags                      BufferCreateFlags
    size                       DeviceSize
    usage                      BufferUsageFlags
    sharing_mode               SharingMode
    queue_family_index_count   u32
    p_queue_family_indices     &u32
} 

pub struct BufferViewCreateInfo {
mut:
    s_type                         StructureType
    p_next                         voidptr
    flags                          BufferViewCreateFlags
    buffer                         C.Buffer
    format                         Format
    offset                         DeviceSize
    range                          DeviceSize
} 

pub struct ImageCreateInfo {
mut:
    s_type                       StructureType
    p_next                       voidptr
    flags                        ImageCreateFlags
    image_type                   ImageType
    format                       Format
    extent                       Extent3D
    mip_levels                   u32
    array_layers                 u32
    samples                      SampleCountFlagBits
    tiling                       ImageTiling
    usage                        ImageUsageFlags
    sharing_mode                 SharingMode
    queue_family_index_count     u32
    p_queue_family_indices       &u32
    initial_layout               ImageLayout
} 

pub struct SubresourceLayout {
mut:
    offset              DeviceSize
    size                DeviceSize
    row_pitch           DeviceSize
    array_pitch         DeviceSize
    depth_pitch         DeviceSize
} 

pub struct ComponentMapping {
mut:
    r                         ComponentSwizzle
    g                         ComponentSwizzle
    b                         ComponentSwizzle
    a                         ComponentSwizzle
} 

pub struct ImageViewCreateInfo {
mut:
    s_type                         StructureType
    p_next                         voidptr
    flags                          ImageViewCreateFlags
    image                          C.Image
    view_type                      ImageViewType
    format                         Format
    components                     ComponentMapping
    subresource_range              ImageSubresourceRange
} 

// ShaderModuleCreateInfo extends VkPipelineShaderStageCreateInfo
pub struct ShaderModuleCreateInfo {
mut:
    s_type                           StructureType
    p_next                           voidptr
    flags                            ShaderModuleCreateFlags
    code_size                        usize
    p_code                           &u32
} 

pub struct PipelineCacheCreateInfo {
mut:
    s_type                            StructureType
    p_next                            voidptr
    flags                             PipelineCacheCreateFlags
    initial_data_size                 usize
    p_initial_data                    voidptr
} 

pub struct SpecializationMapEntry {
mut:
    constant_id     u32
    offset          u32
    size            usize
} 

pub struct SpecializationInfo {
mut:
    map_entry_count                        u32
    p_map_entries                          &SpecializationMapEntry
    data_size                              usize
    p_data                                 voidptr
} 

pub struct PipelineShaderStageCreateInfo {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    flags                                   PipelineShaderStageCreateFlags
    stage                                   ShaderStageFlagBits
    vkmodule                                C.ShaderModule
    p_name                                  &char
    p_specialization_info                   &SpecializationInfo
} 

pub struct ComputePipelineCreateInfo {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    flags                                  PipelineCreateFlags
    stage                                  PipelineShaderStageCreateInfo
    layout                                 C.PipelineLayout
    base_pipeline_handle                   C.Pipeline
    base_pipeline_index                    i32
} 

pub struct VertexInputBindingDescription {
mut:
    binding                  u32
    stride                   u32
    input_rate               VertexInputRate
} 

pub struct VertexInputAttributeDescription {
mut:
    location        u32
    binding         u32
    format          Format
    offset          u32
} 

pub struct PipelineVertexInputStateCreateInfo {
mut:
    s_type                                          StructureType
    p_next                                          voidptr
    flags                                           PipelineVertexInputStateCreateFlags
    vertex_binding_description_count                u32
    p_vertex_binding_descriptions                   &VertexInputBindingDescription
    vertex_attribute_description_count              u32
    p_vertex_attribute_descriptions                 &VertexInputAttributeDescription
} 

pub struct PipelineInputAssemblyStateCreateInfo {
mut:
    s_type                                         StructureType
    p_next                                         voidptr
    flags                                          PipelineInputAssemblyStateCreateFlags
    topology                                       PrimitiveTopology
    primitive_restart_enable                       Bool32
} 

pub struct PipelineTessellationStateCreateInfo {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    flags                                         PipelineTessellationStateCreateFlags
    patch_control_points                          u32
} 

pub struct Viewport {
mut:
    x            f32
    y            f32
    width        f32
    height       f32
    min_depth    f32
    max_depth    f32
} 

pub struct PipelineViewportStateCreateInfo {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    flags                                     PipelineViewportStateCreateFlags
    viewport_count                            u32
    p_viewports                               &Viewport
    scissor_count                             u32
    p_scissors                                &Rect2D
} 

pub struct PipelineRasterizationStateCreateInfo {
mut:
    s_type                                         StructureType
    p_next                                         voidptr
    flags                                          PipelineRasterizationStateCreateFlags
    depth_clamp_enable                             Bool32
    rasterizer_discard_enable                      Bool32
    polygon_mode                                   PolygonMode
    cull_mode                                      CullModeFlags
    front_face                                     FrontFace
    depth_bias_enable                              Bool32
    depth_bias_constant_factor                     f32
    depth_bias_clamp                               f32
    depth_bias_slope_factor                        f32
    line_width                                     f32
} 

pub struct PipelineMultisampleStateCreateInfo {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    flags                                        PipelineMultisampleStateCreateFlags
    rasterization_samples                        SampleCountFlagBits
    sample_shading_enable                        Bool32
    min_sample_shading                           f32
    p_sample_mask                                &SampleMask
    alpha_to_coverage_enable                     Bool32
    alpha_to_one_enable                          Bool32
} 

pub struct StencilOpState {
mut:
    fail_op            StencilOp
    pass_op            StencilOp
    depth_fail_op      StencilOp
    compare_op         CompareOp
    compare_mask       u32
    write_mask         u32
    reference          u32
} 

pub struct PipelineDepthStencilStateCreateInfo {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    flags                                         PipelineDepthStencilStateCreateFlags
    depth_test_enable                             Bool32
    depth_write_enable                            Bool32
    depth_compare_op                              CompareOp
    depth_bounds_test_enable                      Bool32
    stencil_test_enable                           Bool32
    front                                         StencilOpState
    back                                          StencilOpState
    min_depth_bounds                              f32
    max_depth_bounds                              f32
} 

pub struct PipelineColorBlendAttachmentState {
mut:
    blend_enable                 Bool32
    src_color_blend_factor       BlendFactor
    dst_color_blend_factor       BlendFactor
    color_blend_op               BlendOp
    src_alpha_blend_factor       BlendFactor
    dst_alpha_blend_factor       BlendFactor
    alpha_blend_op               BlendOp
    color_write_mask             ColorComponentFlags
} 

pub struct PipelineColorBlendStateCreateInfo {
mut:
    s_type                                            StructureType
    p_next                                            voidptr
    flags                                             PipelineColorBlendStateCreateFlags
    logic_op_enable                                   Bool32
    logic_op                                          LogicOp
    attachment_count                                  u32
    p_attachments                                     &PipelineColorBlendAttachmentState
    blend_constants                                   []f32
} 

pub struct PipelineDynamicStateCreateInfo {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    flags                                    PipelineDynamicStateCreateFlags
    dynamic_state_count                      u32
    p_dynamic_states                         &DynamicState
} 

pub struct GraphicsPipelineCreateInfo {
mut:
    s_type                                               StructureType
    p_next                                               voidptr
    flags                                                PipelineCreateFlags
    stage_count                                          u32
    p_stages                                             &PipelineShaderStageCreateInfo
    p_vertex_input_state                                 &PipelineVertexInputStateCreateInfo
    p_input_assembly_state                               &PipelineInputAssemblyStateCreateInfo
    p_tessellation_state                                 &PipelineTessellationStateCreateInfo
    p_viewport_state                                     &PipelineViewportStateCreateInfo
    p_rasterization_state                                &PipelineRasterizationStateCreateInfo
    p_multisample_state                                  &PipelineMultisampleStateCreateInfo
    p_depth_stencil_state                                &PipelineDepthStencilStateCreateInfo
    p_color_blend_state                                  &PipelineColorBlendStateCreateInfo
    p_dynamic_state                                      &PipelineDynamicStateCreateInfo
    layout                                               C.PipelineLayout
    render_pass                                          C.RenderPass
    subpass                                              u32
    base_pipeline_handle                                 C.Pipeline
    base_pipeline_index                                  i32
} 

pub struct PushConstantRange {
mut:
    stage_flags               ShaderStageFlags
    offset                    u32
    size                      u32
} 

pub struct PipelineLayoutCreateInfo {
mut:
    s_type                              StructureType
    p_next                              voidptr
    flags                               PipelineLayoutCreateFlags
    set_layout_count                    u32
    p_set_layouts                       &C.DescriptorSetLayout
    push_constant_range_count           u32
    p_push_constant_ranges              &PushConstantRange
} 

pub struct SamplerCreateInfo {
mut:
    s_type                      StructureType
    p_next                      voidptr
    flags                       SamplerCreateFlags
    mag_filter                  Filter
    min_filter                  Filter
    mipmap_mode                 SamplerMipmapMode
    address_mode_u              SamplerAddressMode
    address_mode_v              SamplerAddressMode
    address_mode_w              SamplerAddressMode
    mip_lod_bias                f32
    anisotropy_enable           Bool32
    max_anisotropy              f32
    compare_enable              Bool32
    compare_op                  CompareOp
    min_lod                     f32
    max_lod                     f32
    border_color                BorderColor
    unnormalized_coordinates    Bool32
} 

pub struct CopyDescriptorSet {
mut:
    s_type                 StructureType
    p_next                 voidptr
    src_set                C.DescriptorSet
    src_binding            u32
    src_array_element      u32
    dst_set                C.DescriptorSet
    dst_binding            u32
    dst_array_element      u32
    descriptor_count       u32
} 

pub struct DescriptorBufferInfo {
mut:
    buffer              C.Buffer
    offset              DeviceSize
    range               DeviceSize
} 

pub struct DescriptorImageInfo {
mut:
    sampler              C.Sampler
    image_view           C.ImageView
    image_layout         ImageLayout
} 

pub struct DescriptorPoolSize {
mut:
    vktype                  DescriptorType
    descriptor_count        u32
} 

pub struct DescriptorPoolCreateInfo {
mut:
    s_type                             StructureType
    p_next                             voidptr
    flags                              DescriptorPoolCreateFlags
    max_sets                           u32
    pool_size_count                    u32
    p_pool_sizes                       &DescriptorPoolSize
} 

pub struct DescriptorSetAllocateInfo {
mut:
    s_type                              StructureType
    p_next                              voidptr
    descriptor_pool                     C.DescriptorPool
    descriptor_set_count                u32
    p_set_layouts                       &C.DescriptorSetLayout
} 

pub struct DescriptorSetLayoutBinding {
mut:
    binding                   u32
    descriptor_type           DescriptorType
    descriptor_count          u32
    stage_flags               ShaderStageFlags
    p_immutable_samplers      &C.Sampler
} 

pub struct DescriptorSetLayoutCreateInfo {
mut:
    s_type                                     StructureType
    p_next                                     voidptr
    flags                                      DescriptorSetLayoutCreateFlags
    binding_count                              u32
    p_bindings                                 &DescriptorSetLayoutBinding
} 

pub struct WriteDescriptorSet {
mut:
    s_type                               StructureType
    p_next                               voidptr
    dst_set                              C.DescriptorSet
    dst_binding                          u32
    dst_array_element                    u32
    descriptor_count                     u32
    descriptor_type                      DescriptorType
    p_image_info                         &DescriptorImageInfo
    p_buffer_info                        &DescriptorBufferInfo
    p_texel_buffer_view                  &C.BufferView
} 

pub struct AttachmentDescription {
mut:
    flags                               AttachmentDescriptionFlags
    format                              Format
    samples                             SampleCountFlagBits
    load_op                             AttachmentLoadOp
    store_op                            AttachmentStoreOp
    stencil_load_op                     AttachmentLoadOp
    stencil_store_op                    AttachmentStoreOp
    initial_layout                      ImageLayout
    final_layout                        ImageLayout
} 

pub struct AttachmentReference {
mut:
    attachment           u32
    layout               ImageLayout
} 

pub struct FramebufferCreateInfo {
mut:
    s_type                          StructureType
    p_next                          voidptr
    flags                           FramebufferCreateFlags
    render_pass                     C.RenderPass
    attachment_count                u32
    p_attachments                   &C.ImageView
    width                           u32
    height                          u32
    layers                          u32
} 

pub struct SubpassDescription {
mut:
    flags                               SubpassDescriptionFlags
    pipeline_bind_point                 PipelineBindPoint
    input_attachment_count              u32
    p_input_attachments                 &AttachmentReference
    color_attachment_count              u32
    p_color_attachments                 &AttachmentReference
    p_resolve_attachments               &AttachmentReference
    p_depth_stencil_attachment          &AttachmentReference
    preserve_attachment_count           u32
    p_preserve_attachments              &u32
} 

pub struct SubpassDependency {
mut:
    src_subpass                 u32
    dst_subpass                 u32
    src_stage_mask              PipelineStageFlags
    dst_stage_mask              PipelineStageFlags
    src_access_mask             AccessFlags
    dst_access_mask             AccessFlags
    dependency_flags            DependencyFlags
} 

pub struct RenderPassCreateInfo {
mut:
    s_type                                StructureType
    p_next                                voidptr
    flags                                 RenderPassCreateFlags
    attachment_count                      u32
    p_attachments                         &AttachmentDescription
    subpass_count                         u32
    p_subpasses                           &SubpassDescription
    dependency_count                      u32
    p_dependencies                        &SubpassDependency
} 

pub struct CommandPoolCreateInfo {
mut:
    s_type                          StructureType
    p_next                          voidptr
    flags                           CommandPoolCreateFlags
    queue_family_index              u32
} 

pub struct CommandBufferAllocateInfo {
mut:
    s_type                      StructureType
    p_next                      voidptr
    command_pool                C.CommandPool
    level                       CommandBufferLevel
    command_buffer_count        u32
} 

pub struct CommandBufferInheritanceInfo {
mut:
    s_type                               StructureType
    p_next                               voidptr
    render_pass                          C.RenderPass
    subpass                              u32
    framebuffer                          C.Framebuffer
    occlusion_query_enable               Bool32
    query_flags                          QueryControlFlags
    pipeline_statistics                  QueryPipelineStatisticFlags
} 

pub struct CommandBufferBeginInfo {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    flags                                        CommandBufferUsageFlags
    p_inheritance_info                           &CommandBufferInheritanceInfo
} 

pub struct BufferCopy {
mut:
    src_offset          DeviceSize
    dst_offset          DeviceSize
    size                DeviceSize
} 

pub struct ImageSubresourceLayers {
mut:
    aspect_mask               ImageAspectFlags
    mip_level                 u32
    base_array_layer          u32
    layer_count               u32
} 

pub struct BufferImageCopy {
mut:
    buffer_offset                   DeviceSize
    buffer_row_length               u32
    buffer_image_height             u32
    image_subresource               ImageSubresourceLayers
    image_offset                    Offset3D
    image_extent                    Extent3D
} 

pub union ClearColorValue {
mut:
    float32         []f32
    int32           []i32
    uint32          []u32
} 

pub struct ClearDepthStencilValue {
mut:
    depth           f32
    stencil         u32
} 

pub union ClearValue {
mut:
    color                           ClearColorValue
    depth_stencil                   ClearDepthStencilValue
} 

pub struct ClearAttachment {
mut:
    aspect_mask               ImageAspectFlags
    color_attachment          u32
    clear_value               ClearValue
} 

pub struct ClearRect {
mut:
    rect            Rect2D
    base_array_layer u32
    layer_count     u32
} 

pub struct ImageBlit {
mut:
    src_subresource                 ImageSubresourceLayers
    src_offsets                     []Offset3D
    dst_subresource                 ImageSubresourceLayers
    dst_offsets                     []Offset3D
} 

pub struct ImageCopy {
mut:
    src_subresource                 ImageSubresourceLayers
    src_offset                      Offset3D
    dst_subresource                 ImageSubresourceLayers
    dst_offset                      Offset3D
    extent                          Extent3D
} 

pub struct ImageResolve {
mut:
    src_subresource                 ImageSubresourceLayers
    src_offset                      Offset3D
    dst_subresource                 ImageSubresourceLayers
    dst_offset                      Offset3D
    extent                          Extent3D
} 

pub struct RenderPassBeginInfo {
mut:
    s_type                     StructureType
    p_next                     voidptr
    render_pass                C.RenderPass
    framebuffer                C.Framebuffer
    render_area                Rect2D
    clear_value_count          u32
    p_clear_values             &ClearValue
} 

type VkCreateInstance = fn (     &InstanceCreateInfo,     &AllocationCallbacks,     &C.Instance) Result

pub fn create_instance(
    p_create_info                                   &InstanceCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_instance                                      &C.Instance) Result {
      f := VkCreateInstance((*loader_p).get_sym('vkCreateInstance'
    ) or { 
        println("Couldn't load symbol for 'vkCreateInstance': ${err}")
        return Result.error_unknown
    })
    return f(
    p_create_info,
    p_allocator,
    p_instance)
}


type VkDestroyInstance = fn (     C.Instance,     &AllocationCallbacks) 

pub fn destroy_instance(
    instance                                        C.Instance,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyInstance((*loader_p).get_sym('vkDestroyInstance'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyInstance': ${err}")
        return 
    })
    f(
    instance,
    p_allocator)
}


type VkEnumeratePhysicalDevices = fn (     C.Instance,     &u32,     &C.PhysicalDevice) Result

pub fn enumerate_physical_devices(
    instance                                        C.Instance,
    p_physical_device_count                         &u32,
    p_physical_devices                              &C.PhysicalDevice) Result {
      f := VkEnumeratePhysicalDevices((*loader_p).get_sym('vkEnumeratePhysicalDevices'
    ) or { 
        println("Couldn't load symbol for 'vkEnumeratePhysicalDevices': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_physical_device_count,
    p_physical_devices)
}


type VkGetPhysicalDeviceFeatures = fn (     C.PhysicalDevice,     &PhysicalDeviceFeatures) 

pub fn get_physical_device_features(
    physical_device                                 C.PhysicalDevice,
    p_features                                      &PhysicalDeviceFeatures)  {
      f := VkGetPhysicalDeviceFeatures((*loader_p).get_sym('vkGetPhysicalDeviceFeatures'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceFeatures': ${err}")
        return 
    })
    f(
    physical_device,
    p_features)
}


type VkGetPhysicalDeviceFormatProperties = fn (     C.PhysicalDevice,     Format,     &FormatProperties) 

pub fn get_physical_device_format_properties(
    physical_device                                 C.PhysicalDevice,
    format                                          Format,
    p_format_properties                             &FormatProperties)  {
      f := VkGetPhysicalDeviceFormatProperties((*loader_p).get_sym('vkGetPhysicalDeviceFormatProperties'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceFormatProperties': ${err}")
        return 
    })
    f(
    physical_device,
    format,
    p_format_properties)
}


type VkGetPhysicalDeviceImageFormatProperties = fn (     C.PhysicalDevice,     Format,     ImageType,     ImageTiling,     ImageUsageFlags,     ImageCreateFlags,     &ImageFormatProperties) Result

pub fn get_physical_device_image_format_properties(
    physical_device                                 C.PhysicalDevice,
    format                                          Format,
    vktype                                          ImageType,
    tiling                                          ImageTiling,
    usage                                           ImageUsageFlags,
    flags                                           ImageCreateFlags,
    p_image_format_properties                       &ImageFormatProperties) Result {
      f := VkGetPhysicalDeviceImageFormatProperties((*loader_p).get_sym('vkGetPhysicalDeviceImageFormatProperties'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceImageFormatProperties': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    format,
    vktype,
    tiling,
    usage,
    flags,
    p_image_format_properties)
}


type VkGetPhysicalDeviceProperties = fn (     C.PhysicalDevice,     &PhysicalDeviceProperties) 

pub fn get_physical_device_properties(
    physical_device                                 C.PhysicalDevice,
    p_properties                                    &PhysicalDeviceProperties)  {
      f := VkGetPhysicalDeviceProperties((*loader_p).get_sym('vkGetPhysicalDeviceProperties'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceProperties': ${err}")
        return 
    })
    f(
    physical_device,
    p_properties)
}


type VkGetPhysicalDeviceQueueFamilyProperties = fn (     C.PhysicalDevice,     &u32,     &QueueFamilyProperties) 

pub fn get_physical_device_queue_family_properties(
    physical_device                                 C.PhysicalDevice,
    p_queue_family_property_count                   &u32,
    p_queue_family_properties                       &QueueFamilyProperties)  {
      f := VkGetPhysicalDeviceQueueFamilyProperties((*loader_p).get_sym('vkGetPhysicalDeviceQueueFamilyProperties'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceQueueFamilyProperties': ${err}")
        return 
    })
    f(
    physical_device,
    p_queue_family_property_count,
    p_queue_family_properties)
}


type VkGetPhysicalDeviceMemoryProperties = fn (     C.PhysicalDevice,     &PhysicalDeviceMemoryProperties) 

pub fn get_physical_device_memory_properties(
    physical_device                                 C.PhysicalDevice,
    p_memory_properties                             &PhysicalDeviceMemoryProperties)  {
      f := VkGetPhysicalDeviceMemoryProperties((*loader_p).get_sym('vkGetPhysicalDeviceMemoryProperties'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceMemoryProperties': ${err}")
        return 
    })
    f(
    physical_device,
    p_memory_properties)
}


type VkGetInstanceProcAddr = fn (     C.Instance,     &char) PFN_vkVoidFunction

pub fn get_instance_proc_addr(
    instance                                        C.Instance,
    p_name                                          &char) PFN_vkVoidFunction {
      f := VkGetInstanceProcAddr((*loader_p).get_sym("vkGetInstanceProcAddr"
    ) or { 
        panic("Couldn't load symbol for 'vkGetInstanceProcAddr': ${err}") })
    return f(
    instance,
    p_name)
}


type VkGetDeviceProcAddr = fn (     C.Device,     &char) PFN_vkVoidFunction

pub fn get_device_proc_addr(
    device                                          C.Device,
    p_name                                          &char) PFN_vkVoidFunction {
      f := VkGetDeviceProcAddr((*loader_p).get_sym("vkGetDeviceProcAddr"
    ) or { 
        panic("Couldn't load symbol for 'vkGetDeviceProcAddr': ${err}") })
    return f(
    device,
    p_name)
}


type VkCreateDevice = fn (     C.PhysicalDevice,     &DeviceCreateInfo,     &AllocationCallbacks,     &C.Device) Result

pub fn create_device(
    physical_device                                 C.PhysicalDevice,
    p_create_info                                   &DeviceCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_device                                        &C.Device) Result {
      f := VkCreateDevice((*loader_p).get_sym('vkCreateDevice'
    ) or { 
        println("Couldn't load symbol for 'vkCreateDevice': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_create_info,
    p_allocator,
    p_device)
}


type VkDestroyDevice = fn (     C.Device,     &AllocationCallbacks) 

pub fn destroy_device(
    device                                          C.Device,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyDevice((*loader_p).get_sym('vkDestroyDevice'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyDevice': ${err}")
        return 
    })
    f(
    device,
    p_allocator)
}


type VkEnumerateInstanceExtensionProperties = fn (     &char,     &u32,     &ExtensionProperties) Result

pub fn enumerate_instance_extension_properties(
    p_layer_name                                    &char,
    p_property_count                                &u32,
    p_properties                                    &ExtensionProperties) Result {
      f := VkEnumerateInstanceExtensionProperties((*loader_p).get_sym('vkEnumerateInstanceExtensionProperties'
    ) or { 
        println("Couldn't load symbol for 'vkEnumerateInstanceExtensionProperties': ${err}")
        return Result.error_unknown
    })
    return f(
    p_layer_name,
    p_property_count,
    p_properties)
}


type VkEnumerateDeviceExtensionProperties = fn (     C.PhysicalDevice,     &char,     &u32,     &ExtensionProperties) Result

pub fn enumerate_device_extension_properties(
    physical_device                                 C.PhysicalDevice,
    p_layer_name                                    &char,
    p_property_count                                &u32,
    p_properties                                    &ExtensionProperties) Result {
      f := VkEnumerateDeviceExtensionProperties((*loader_p).get_sym('vkEnumerateDeviceExtensionProperties'
    ) or { 
        println("Couldn't load symbol for 'vkEnumerateDeviceExtensionProperties': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_layer_name,
    p_property_count,
    p_properties)
}


type VkEnumerateInstanceLayerProperties = fn (     &u32,     &LayerProperties) Result

pub fn enumerate_instance_layer_properties(
    p_property_count                                &u32,
    p_properties                                    &LayerProperties) Result {
      f := VkEnumerateInstanceLayerProperties((*loader_p).get_sym('vkEnumerateInstanceLayerProperties'
    ) or { 
        println("Couldn't load symbol for 'vkEnumerateInstanceLayerProperties': ${err}")
        return Result.error_unknown
    })
    return f(
    p_property_count,
    p_properties)
}


type VkEnumerateDeviceLayerProperties = fn (     C.PhysicalDevice,     &u32,     &LayerProperties) Result

pub fn enumerate_device_layer_properties(
    physical_device                                 C.PhysicalDevice,
    p_property_count                                &u32,
    p_properties                                    &LayerProperties) Result {
      f := VkEnumerateDeviceLayerProperties((*loader_p).get_sym('vkEnumerateDeviceLayerProperties'
    ) or { 
        println("Couldn't load symbol for 'vkEnumerateDeviceLayerProperties': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_property_count,
    p_properties)
}


type VkGetDeviceQueue = fn (     C.Device,     u32,     u32,     &C.Queue) 

pub fn get_device_queue(
    device                                          C.Device,
    queue_family_index                              u32,
    queue_index                                     u32,
    p_queue                                         &C.Queue)  {
      f := VkGetDeviceQueue((*loader_p).get_sym('vkGetDeviceQueue'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceQueue': ${err}")
        return 
    })
    f(
    device,
    queue_family_index,
    queue_index,
    p_queue)
}


type VkQueueSubmit = fn (     C.Queue,     u32,     &SubmitInfo,     C.Fence) Result

pub fn queue_submit(
    queue                                           C.Queue,
    submit_count                                    u32,
    p_submits                                       &SubmitInfo,
    fence                                           C.Fence) Result {
      f := VkQueueSubmit((*loader_p).get_sym('vkQueueSubmit'
    ) or { 
        println("Couldn't load symbol for 'vkQueueSubmit': ${err}")
        return Result.error_unknown
    })
    return f(
    queue,
    submit_count,
    p_submits,
    fence)
}


type VkQueueWaitIdle = fn (     C.Queue) Result

pub fn queue_wait_idle(
    queue                                           C.Queue) Result {
      f := VkQueueWaitIdle((*loader_p).get_sym('vkQueueWaitIdle'
    ) or { 
        println("Couldn't load symbol for 'vkQueueWaitIdle': ${err}")
        return Result.error_unknown
    })
    return f(
    queue)
}


type VkDeviceWaitIdle = fn (     C.Device) Result

pub fn device_wait_idle(
    device                                          C.Device) Result {
      f := VkDeviceWaitIdle((*loader_p).get_sym('vkDeviceWaitIdle'
    ) or { 
        println("Couldn't load symbol for 'vkDeviceWaitIdle': ${err}")
        return Result.error_unknown
    })
    return f(
    device)
}


type VkAllocateMemory = fn (     C.Device,     &MemoryAllocateInfo,     &AllocationCallbacks,     &C.DeviceMemory) Result

pub fn allocate_memory(
    device                                          C.Device,
    p_allocate_info                                 &MemoryAllocateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_memory                                        &C.DeviceMemory) Result {
      f := VkAllocateMemory((*loader_p).get_sym('vkAllocateMemory'
    ) or { 
        println("Couldn't load symbol for 'vkAllocateMemory': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_allocate_info,
    p_allocator,
    p_memory)
}


type VkFreeMemory = fn (     C.Device,     C.DeviceMemory,     &AllocationCallbacks) 

pub fn free_memory(
    device                                          C.Device,
    memory                                          C.DeviceMemory,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkFreeMemory((*loader_p).get_sym('vkFreeMemory'
    ) or { 
        println("Couldn't load symbol for 'vkFreeMemory': ${err}")
        return 
    })
    f(
    device,
    memory,
    p_allocator)
}


type VkMapMemory = fn (     C.Device,     C.DeviceMemory,     DeviceSize,     DeviceSize,     MemoryMapFlags,     &voidptr) Result

pub fn map_memory(
    device                                          C.Device,
    memory                                          C.DeviceMemory,
    offset                                          DeviceSize,
    size                                            DeviceSize,
    flags                                           MemoryMapFlags,
    pp_data                                         &voidptr) Result {
      f := VkMapMemory((*loader_p).get_sym('vkMapMemory'
    ) or { 
        println("Couldn't load symbol for 'vkMapMemory': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    memory,
    offset,
    size,
    flags,
    pp_data)
}


type VkUnmapMemory = fn (     C.Device,     C.DeviceMemory) 

pub fn unmap_memory(
    device                                          C.Device,
    memory                                          C.DeviceMemory)  {
      f := VkUnmapMemory((*loader_p).get_sym('vkUnmapMemory'
    ) or { 
        println("Couldn't load symbol for 'vkUnmapMemory': ${err}")
        return 
    })
    f(
    device,
    memory)
}


type VkFlushMappedMemoryRanges = fn (     C.Device,     u32,     &MappedMemoryRange) Result

pub fn flush_mapped_memory_ranges(
    device                                          C.Device,
    memory_range_count                              u32,
    p_memory_ranges                                 &MappedMemoryRange) Result {
      f := VkFlushMappedMemoryRanges((*loader_p).get_sym('vkFlushMappedMemoryRanges'
    ) or { 
        println("Couldn't load symbol for 'vkFlushMappedMemoryRanges': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    memory_range_count,
    p_memory_ranges)
}


type VkInvalidateMappedMemoryRanges = fn (     C.Device,     u32,     &MappedMemoryRange) Result

pub fn invalidate_mapped_memory_ranges(
    device                                          C.Device,
    memory_range_count                              u32,
    p_memory_ranges                                 &MappedMemoryRange) Result {
      f := VkInvalidateMappedMemoryRanges((*loader_p).get_sym('vkInvalidateMappedMemoryRanges'
    ) or { 
        println("Couldn't load symbol for 'vkInvalidateMappedMemoryRanges': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    memory_range_count,
    p_memory_ranges)
}


type VkGetDeviceMemoryCommitment = fn (     C.Device,     C.DeviceMemory,     &DeviceSize) 

pub fn get_device_memory_commitment(
    device                                          C.Device,
    memory                                          C.DeviceMemory,
    p_committed_memory_in_bytes                     &DeviceSize)  {
      f := VkGetDeviceMemoryCommitment((*loader_p).get_sym('vkGetDeviceMemoryCommitment'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceMemoryCommitment': ${err}")
        return 
    })
    f(
    device,
    memory,
    p_committed_memory_in_bytes)
}


type VkBindBufferMemory = fn (     C.Device,     C.Buffer,     C.DeviceMemory,     DeviceSize) Result

pub fn bind_buffer_memory(
    device                                          C.Device,
    buffer                                          C.Buffer,
    memory                                          C.DeviceMemory,
    memory_offset                                   DeviceSize) Result {
      f := VkBindBufferMemory((*loader_p).get_sym('vkBindBufferMemory'
    ) or { 
        println("Couldn't load symbol for 'vkBindBufferMemory': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    buffer,
    memory,
    memory_offset)
}


type VkBindImageMemory = fn (     C.Device,     C.Image,     C.DeviceMemory,     DeviceSize) Result

pub fn bind_image_memory(
    device                                          C.Device,
    image                                           C.Image,
    memory                                          C.DeviceMemory,
    memory_offset                                   DeviceSize) Result {
      f := VkBindImageMemory((*loader_p).get_sym('vkBindImageMemory'
    ) or { 
        println("Couldn't load symbol for 'vkBindImageMemory': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    image,
    memory,
    memory_offset)
}


type VkGetBufferMemoryRequirements = fn (     C.Device,     C.Buffer,     &MemoryRequirements) 

pub fn get_buffer_memory_requirements(
    device                                          C.Device,
    buffer                                          C.Buffer,
    p_memory_requirements                           &MemoryRequirements)  {
      f := VkGetBufferMemoryRequirements((*loader_p).get_sym('vkGetBufferMemoryRequirements'
    ) or { 
        println("Couldn't load symbol for 'vkGetBufferMemoryRequirements': ${err}")
        return 
    })
    f(
    device,
    buffer,
    p_memory_requirements)
}


type VkGetImageMemoryRequirements = fn (     C.Device,     C.Image,     &MemoryRequirements) 

pub fn get_image_memory_requirements(
    device                                          C.Device,
    image                                           C.Image,
    p_memory_requirements                           &MemoryRequirements)  {
      f := VkGetImageMemoryRequirements((*loader_p).get_sym('vkGetImageMemoryRequirements'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageMemoryRequirements': ${err}")
        return 
    })
    f(
    device,
    image,
    p_memory_requirements)
}


type VkGetImageSparseMemoryRequirements = fn (     C.Device,     C.Image,     &u32,     &SparseImageMemoryRequirements) 

pub fn get_image_sparse_memory_requirements(
    device                                          C.Device,
    image                                           C.Image,
    p_sparse_memory_requirement_count               &u32,
    p_sparse_memory_requirements                    &SparseImageMemoryRequirements)  {
      f := VkGetImageSparseMemoryRequirements((*loader_p).get_sym('vkGetImageSparseMemoryRequirements'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageSparseMemoryRequirements': ${err}")
        return 
    })
    f(
    device,
    image,
    p_sparse_memory_requirement_count,
    p_sparse_memory_requirements)
}


type VkGetPhysicalDeviceSparseImageFormatProperties = fn (     C.PhysicalDevice,     Format,     ImageType,     SampleCountFlagBits,     ImageUsageFlags,     ImageTiling,     &u32,     &SparseImageFormatProperties) 

pub fn get_physical_device_sparse_image_format_properties(
    physical_device                                 C.PhysicalDevice,
    format                                          Format,
    vktype                                          ImageType,
    samples                                         SampleCountFlagBits,
    usage                                           ImageUsageFlags,
    tiling                                          ImageTiling,
    p_property_count                                &u32,
    p_properties                                    &SparseImageFormatProperties)  {
      f := VkGetPhysicalDeviceSparseImageFormatProperties((*loader_p).get_sym('vkGetPhysicalDeviceSparseImageFormatProperties'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSparseImageFormatProperties': ${err}")
        return 
    })
    f(
    physical_device,
    format,
    vktype,
    samples,
    usage,
    tiling,
    p_property_count,
    p_properties)
}


type VkQueueBindSparse = fn (     C.Queue,     u32,     &BindSparseInfo,     C.Fence) Result

pub fn queue_bind_sparse(
    queue                                           C.Queue,
    bind_info_count                                 u32,
    p_bind_info                                     &BindSparseInfo,
    fence                                           C.Fence) Result {
      f := VkQueueBindSparse((*loader_p).get_sym('vkQueueBindSparse'
    ) or { 
        println("Couldn't load symbol for 'vkQueueBindSparse': ${err}")
        return Result.error_unknown
    })
    return f(
    queue,
    bind_info_count,
    p_bind_info,
    fence)
}


type VkCreateFence = fn (     C.Device,     &FenceCreateInfo,     &AllocationCallbacks,     &C.Fence) Result

pub fn create_fence(
    device                                          C.Device,
    p_create_info                                   &FenceCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_fence                                         &C.Fence) Result {
      f := VkCreateFence((*loader_p).get_sym('vkCreateFence'
    ) or { 
        println("Couldn't load symbol for 'vkCreateFence': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_fence)
}


type VkDestroyFence = fn (     C.Device,     C.Fence,     &AllocationCallbacks) 

pub fn destroy_fence(
    device                                          C.Device,
    fence                                           C.Fence,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyFence((*loader_p).get_sym('vkDestroyFence'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyFence': ${err}")
        return 
    })
    f(
    device,
    fence,
    p_allocator)
}


type VkResetFences = fn (     C.Device,     u32,     &C.Fence) Result

pub fn reset_fences(
    device                                          C.Device,
    fence_count                                     u32,
    p_fences                                        &C.Fence) Result {
      f := VkResetFences((*loader_p).get_sym('vkResetFences'
    ) or { 
        println("Couldn't load symbol for 'vkResetFences': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    fence_count,
    p_fences)
}


type VkGetFenceStatus = fn (     C.Device,     C.Fence) Result

pub fn get_fence_status(
    device                                          C.Device,
    fence                                           C.Fence) Result {
      f := VkGetFenceStatus((*loader_p).get_sym('vkGetFenceStatus'
    ) or { 
        println("Couldn't load symbol for 'vkGetFenceStatus': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    fence)
}


type VkWaitForFences = fn (     C.Device,     u32,     &C.Fence,     Bool32,     u64) Result

pub fn wait_for_fences(
    device                                          C.Device,
    fence_count                                     u32,
    p_fences                                        &C.Fence,
    wait_all                                        Bool32,
    timeout                                         u64) Result {
      f := VkWaitForFences((*loader_p).get_sym('vkWaitForFences'
    ) or { 
        println("Couldn't load symbol for 'vkWaitForFences': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    fence_count,
    p_fences,
    wait_all,
    timeout)
}


type VkCreateSemaphore = fn (     C.Device,     &SemaphoreCreateInfo,     &AllocationCallbacks,     &C.Semaphore) Result

pub fn create_semaphore(
    device                                          C.Device,
    p_create_info                                   &SemaphoreCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_semaphore                                     &C.Semaphore) Result {
      f := VkCreateSemaphore((*loader_p).get_sym('vkCreateSemaphore'
    ) or { 
        println("Couldn't load symbol for 'vkCreateSemaphore': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_semaphore)
}


type VkDestroySemaphore = fn (     C.Device,     C.Semaphore,     &AllocationCallbacks) 

pub fn destroy_semaphore(
    device                                          C.Device,
    semaphore                                       C.Semaphore,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroySemaphore((*loader_p).get_sym('vkDestroySemaphore'
    ) or { 
        println("Couldn't load symbol for 'vkDestroySemaphore': ${err}")
        return 
    })
    f(
    device,
    semaphore,
    p_allocator)
}


type VkCreateEvent = fn (     C.Device,     &EventCreateInfo,     &AllocationCallbacks,     &C.Event) Result

pub fn create_event(
    device                                          C.Device,
    p_create_info                                   &EventCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_event                                         &C.Event) Result {
      f := VkCreateEvent((*loader_p).get_sym('vkCreateEvent'
    ) or { 
        println("Couldn't load symbol for 'vkCreateEvent': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_event)
}


type VkDestroyEvent = fn (     C.Device,     C.Event,     &AllocationCallbacks) 

pub fn destroy_event(
    device                                          C.Device,
    event                                           C.Event,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyEvent((*loader_p).get_sym('vkDestroyEvent'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyEvent': ${err}")
        return 
    })
    f(
    device,
    event,
    p_allocator)
}


type VkGetEventStatus = fn (     C.Device,     C.Event) Result

pub fn get_event_status(
    device                                          C.Device,
    event                                           C.Event) Result {
      f := VkGetEventStatus((*loader_p).get_sym('vkGetEventStatus'
    ) or { 
        println("Couldn't load symbol for 'vkGetEventStatus': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    event)
}


type VkSetEvent = fn (     C.Device,     C.Event) Result

pub fn set_event(
    device                                          C.Device,
    event                                           C.Event) Result {
      f := VkSetEvent((*loader_p).get_sym('vkSetEvent'
    ) or { 
        println("Couldn't load symbol for 'vkSetEvent': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    event)
}


type VkResetEvent = fn (     C.Device,     C.Event) Result

pub fn reset_event(
    device                                          C.Device,
    event                                           C.Event) Result {
      f := VkResetEvent((*loader_p).get_sym('vkResetEvent'
    ) or { 
        println("Couldn't load symbol for 'vkResetEvent': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    event)
}


type VkCreateQueryPool = fn (     C.Device,     &QueryPoolCreateInfo,     &AllocationCallbacks,     &C.QueryPool) Result

pub fn create_query_pool(
    device                                          C.Device,
    p_create_info                                   &QueryPoolCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_query_pool                                    &C.QueryPool) Result {
      f := VkCreateQueryPool((*loader_p).get_sym('vkCreateQueryPool'
    ) or { 
        println("Couldn't load symbol for 'vkCreateQueryPool': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_query_pool)
}


type VkDestroyQueryPool = fn (     C.Device,     C.QueryPool,     &AllocationCallbacks) 

pub fn destroy_query_pool(
    device                                          C.Device,
    query_pool                                      C.QueryPool,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyQueryPool((*loader_p).get_sym('vkDestroyQueryPool'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyQueryPool': ${err}")
        return 
    })
    f(
    device,
    query_pool,
    p_allocator)
}


type VkGetQueryPoolResults = fn (     C.Device,     C.QueryPool,     u32,     u32,     usize,     voidptr,     DeviceSize,     QueryResultFlags) Result

pub fn get_query_pool_results(
    device                                          C.Device,
    query_pool                                      C.QueryPool,
    first_query                                     u32,
    query_count                                     u32,
    data_size                                       usize,
    p_data                                          voidptr,
    stride                                          DeviceSize,
    flags                                           QueryResultFlags) Result {
      f := VkGetQueryPoolResults((*loader_p).get_sym('vkGetQueryPoolResults'
    ) or { 
        println("Couldn't load symbol for 'vkGetQueryPoolResults': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    query_pool,
    first_query,
    query_count,
    data_size,
    p_data,
    stride,
    flags)
}


type VkCreateBuffer = fn (     C.Device,     &BufferCreateInfo,     &AllocationCallbacks,     &C.Buffer) Result

pub fn create_buffer(
    device                                          C.Device,
    p_create_info                                   &BufferCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_buffer                                        &C.Buffer) Result {
      f := VkCreateBuffer((*loader_p).get_sym('vkCreateBuffer'
    ) or { 
        println("Couldn't load symbol for 'vkCreateBuffer': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_buffer)
}


type VkDestroyBuffer = fn (     C.Device,     C.Buffer,     &AllocationCallbacks) 

pub fn destroy_buffer(
    device                                          C.Device,
    buffer                                          C.Buffer,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyBuffer((*loader_p).get_sym('vkDestroyBuffer'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyBuffer': ${err}")
        return 
    })
    f(
    device,
    buffer,
    p_allocator)
}


type VkCreateBufferView = fn (     C.Device,     &BufferViewCreateInfo,     &AllocationCallbacks,     &C.BufferView) Result

pub fn create_buffer_view(
    device                                          C.Device,
    p_create_info                                   &BufferViewCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_view                                          &C.BufferView) Result {
      f := VkCreateBufferView((*loader_p).get_sym('vkCreateBufferView'
    ) or { 
        println("Couldn't load symbol for 'vkCreateBufferView': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_view)
}


type VkDestroyBufferView = fn (     C.Device,     C.BufferView,     &AllocationCallbacks) 

pub fn destroy_buffer_view(
    device                                          C.Device,
    buffer_view                                     C.BufferView,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyBufferView((*loader_p).get_sym('vkDestroyBufferView'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyBufferView': ${err}")
        return 
    })
    f(
    device,
    buffer_view,
    p_allocator)
}


type VkCreateImage = fn (     C.Device,     &ImageCreateInfo,     &AllocationCallbacks,     &C.Image) Result

pub fn create_image(
    device                                          C.Device,
    p_create_info                                   &ImageCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_image                                         &C.Image) Result {
      f := VkCreateImage((*loader_p).get_sym('vkCreateImage'
    ) or { 
        println("Couldn't load symbol for 'vkCreateImage': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_image)
}


type VkDestroyImage = fn (     C.Device,     C.Image,     &AllocationCallbacks) 

pub fn destroy_image(
    device                                          C.Device,
    image                                           C.Image,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyImage((*loader_p).get_sym('vkDestroyImage'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyImage': ${err}")
        return 
    })
    f(
    device,
    image,
    p_allocator)
}


type VkGetImageSubresourceLayout = fn (     C.Device,     C.Image,     &ImageSubresource,     &SubresourceLayout) 

pub fn get_image_subresource_layout(
    device                                          C.Device,
    image                                           C.Image,
    p_subresource                                   &ImageSubresource,
    p_layout                                        &SubresourceLayout)  {
      f := VkGetImageSubresourceLayout((*loader_p).get_sym('vkGetImageSubresourceLayout'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageSubresourceLayout': ${err}")
        return 
    })
    f(
    device,
    image,
    p_subresource,
    p_layout)
}


type VkCreateImageView = fn (     C.Device,     &ImageViewCreateInfo,     &AllocationCallbacks,     &C.ImageView) Result

pub fn create_image_view(
    device                                          C.Device,
    p_create_info                                   &ImageViewCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_view                                          &C.ImageView) Result {
      f := VkCreateImageView((*loader_p).get_sym('vkCreateImageView'
    ) or { 
        println("Couldn't load symbol for 'vkCreateImageView': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_view)
}


type VkDestroyImageView = fn (     C.Device,     C.ImageView,     &AllocationCallbacks) 

pub fn destroy_image_view(
    device                                          C.Device,
    image_view                                      C.ImageView,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyImageView((*loader_p).get_sym('vkDestroyImageView'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyImageView': ${err}")
        return 
    })
    f(
    device,
    image_view,
    p_allocator)
}


type VkCreateShaderModule = fn (     C.Device,     &ShaderModuleCreateInfo,     &AllocationCallbacks,     &C.ShaderModule) Result

pub fn create_shader_module(
    device                                          C.Device,
    p_create_info                                   &ShaderModuleCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_shader_module                                 &C.ShaderModule) Result {
      f := VkCreateShaderModule((*loader_p).get_sym('vkCreateShaderModule'
    ) or { 
        println("Couldn't load symbol for 'vkCreateShaderModule': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_shader_module)
}


type VkDestroyShaderModule = fn (     C.Device,     C.ShaderModule,     &AllocationCallbacks) 

pub fn destroy_shader_module(
    device                                          C.Device,
    shader_module                                   C.ShaderModule,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyShaderModule((*loader_p).get_sym('vkDestroyShaderModule'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyShaderModule': ${err}")
        return 
    })
    f(
    device,
    shader_module,
    p_allocator)
}


type VkCreatePipelineCache = fn (     C.Device,     &PipelineCacheCreateInfo,     &AllocationCallbacks,     &C.PipelineCache) Result

pub fn create_pipeline_cache(
    device                                          C.Device,
    p_create_info                                   &PipelineCacheCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_pipeline_cache                                &C.PipelineCache) Result {
      f := VkCreatePipelineCache((*loader_p).get_sym('vkCreatePipelineCache'
    ) or { 
        println("Couldn't load symbol for 'vkCreatePipelineCache': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_pipeline_cache)
}


type VkDestroyPipelineCache = fn (     C.Device,     C.PipelineCache,     &AllocationCallbacks) 

pub fn destroy_pipeline_cache(
    device                                          C.Device,
    pipeline_cache                                  C.PipelineCache,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyPipelineCache((*loader_p).get_sym('vkDestroyPipelineCache'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyPipelineCache': ${err}")
        return 
    })
    f(
    device,
    pipeline_cache,
    p_allocator)
}


type VkGetPipelineCacheData = fn (     C.Device,     C.PipelineCache,     &usize,     voidptr) Result

pub fn get_pipeline_cache_data(
    device                                          C.Device,
    pipeline_cache                                  C.PipelineCache,
    p_data_size                                     &usize,
    p_data                                          voidptr) Result {
      f := VkGetPipelineCacheData((*loader_p).get_sym('vkGetPipelineCacheData'
    ) or { 
        println("Couldn't load symbol for 'vkGetPipelineCacheData': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    pipeline_cache,
    p_data_size,
    p_data)
}


type VkMergePipelineCaches = fn (     C.Device,     C.PipelineCache,     u32,     &C.PipelineCache) Result

pub fn merge_pipeline_caches(
    device                                          C.Device,
    dst_cache                                       C.PipelineCache,
    src_cache_count                                 u32,
    p_src_caches                                    &C.PipelineCache) Result {
      f := VkMergePipelineCaches((*loader_p).get_sym('vkMergePipelineCaches'
    ) or { 
        println("Couldn't load symbol for 'vkMergePipelineCaches': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    dst_cache,
    src_cache_count,
    p_src_caches)
}


type VkCreateGraphicsPipelines = fn (     C.Device,     C.PipelineCache,     u32,     &GraphicsPipelineCreateInfo,     &AllocationCallbacks,     &C.Pipeline) Result

pub fn create_graphics_pipelines(
    device                                          C.Device,
    pipeline_cache                                  C.PipelineCache,
    create_info_count                               u32,
    p_create_infos                                  &GraphicsPipelineCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_pipelines                                     &C.Pipeline) Result {
      f := VkCreateGraphicsPipelines((*loader_p).get_sym('vkCreateGraphicsPipelines'
    ) or { 
        println("Couldn't load symbol for 'vkCreateGraphicsPipelines': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    pipeline_cache,
    create_info_count,
    p_create_infos,
    p_allocator,
    p_pipelines)
}


type VkCreateComputePipelines = fn (     C.Device,     C.PipelineCache,     u32,     &ComputePipelineCreateInfo,     &AllocationCallbacks,     &C.Pipeline) Result

pub fn create_compute_pipelines(
    device                                          C.Device,
    pipeline_cache                                  C.PipelineCache,
    create_info_count                               u32,
    p_create_infos                                  &ComputePipelineCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_pipelines                                     &C.Pipeline) Result {
      f := VkCreateComputePipelines((*loader_p).get_sym('vkCreateComputePipelines'
    ) or { 
        println("Couldn't load symbol for 'vkCreateComputePipelines': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    pipeline_cache,
    create_info_count,
    p_create_infos,
    p_allocator,
    p_pipelines)
}


type VkDestroyPipeline = fn (     C.Device,     C.Pipeline,     &AllocationCallbacks) 

pub fn destroy_pipeline(
    device                                          C.Device,
    pipeline                                        C.Pipeline,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyPipeline((*loader_p).get_sym('vkDestroyPipeline'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyPipeline': ${err}")
        return 
    })
    f(
    device,
    pipeline,
    p_allocator)
}


type VkCreatePipelineLayout = fn (     C.Device,     &PipelineLayoutCreateInfo,     &AllocationCallbacks,     &C.PipelineLayout) Result

pub fn create_pipeline_layout(
    device                                          C.Device,
    p_create_info                                   &PipelineLayoutCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_pipeline_layout                               &C.PipelineLayout) Result {
      f := VkCreatePipelineLayout((*loader_p).get_sym('vkCreatePipelineLayout'
    ) or { 
        println("Couldn't load symbol for 'vkCreatePipelineLayout': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_pipeline_layout)
}


type VkDestroyPipelineLayout = fn (     C.Device,     C.PipelineLayout,     &AllocationCallbacks) 

pub fn destroy_pipeline_layout(
    device                                          C.Device,
    pipeline_layout                                 C.PipelineLayout,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyPipelineLayout((*loader_p).get_sym('vkDestroyPipelineLayout'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyPipelineLayout': ${err}")
        return 
    })
    f(
    device,
    pipeline_layout,
    p_allocator)
}


type VkCreateSampler = fn (     C.Device,     &SamplerCreateInfo,     &AllocationCallbacks,     &C.Sampler) Result

pub fn create_sampler(
    device                                          C.Device,
    p_create_info                                   &SamplerCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_sampler                                       &C.Sampler) Result {
      f := VkCreateSampler((*loader_p).get_sym('vkCreateSampler'
    ) or { 
        println("Couldn't load symbol for 'vkCreateSampler': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_sampler)
}


type VkDestroySampler = fn (     C.Device,     C.Sampler,     &AllocationCallbacks) 

pub fn destroy_sampler(
    device                                          C.Device,
    sampler                                         C.Sampler,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroySampler((*loader_p).get_sym('vkDestroySampler'
    ) or { 
        println("Couldn't load symbol for 'vkDestroySampler': ${err}")
        return 
    })
    f(
    device,
    sampler,
    p_allocator)
}


type VkCreateDescriptorSetLayout = fn (     C.Device,     &DescriptorSetLayoutCreateInfo,     &AllocationCallbacks,     &C.DescriptorSetLayout) Result

pub fn create_descriptor_set_layout(
    device                                          C.Device,
    p_create_info                                   &DescriptorSetLayoutCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_set_layout                                    &C.DescriptorSetLayout) Result {
      f := VkCreateDescriptorSetLayout((*loader_p).get_sym('vkCreateDescriptorSetLayout'
    ) or { 
        println("Couldn't load symbol for 'vkCreateDescriptorSetLayout': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_set_layout)
}


type VkDestroyDescriptorSetLayout = fn (     C.Device,     C.DescriptorSetLayout,     &AllocationCallbacks) 

pub fn destroy_descriptor_set_layout(
    device                                          C.Device,
    descriptor_set_layout                           C.DescriptorSetLayout,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyDescriptorSetLayout((*loader_p).get_sym('vkDestroyDescriptorSetLayout'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyDescriptorSetLayout': ${err}")
        return 
    })
    f(
    device,
    descriptor_set_layout,
    p_allocator)
}


type VkCreateDescriptorPool = fn (     C.Device,     &DescriptorPoolCreateInfo,     &AllocationCallbacks,     &C.DescriptorPool) Result

pub fn create_descriptor_pool(
    device                                          C.Device,
    p_create_info                                   &DescriptorPoolCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_descriptor_pool                               &C.DescriptorPool) Result {
      f := VkCreateDescriptorPool((*loader_p).get_sym('vkCreateDescriptorPool'
    ) or { 
        println("Couldn't load symbol for 'vkCreateDescriptorPool': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_descriptor_pool)
}


type VkDestroyDescriptorPool = fn (     C.Device,     C.DescriptorPool,     &AllocationCallbacks) 

pub fn destroy_descriptor_pool(
    device                                          C.Device,
    descriptor_pool                                 C.DescriptorPool,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyDescriptorPool((*loader_p).get_sym('vkDestroyDescriptorPool'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyDescriptorPool': ${err}")
        return 
    })
    f(
    device,
    descriptor_pool,
    p_allocator)
}


type VkResetDescriptorPool = fn (     C.Device,     C.DescriptorPool,     DescriptorPoolResetFlags) Result

pub fn reset_descriptor_pool(
    device                                          C.Device,
    descriptor_pool                                 C.DescriptorPool,
    flags                                           DescriptorPoolResetFlags) Result {
      f := VkResetDescriptorPool((*loader_p).get_sym('vkResetDescriptorPool'
    ) or { 
        println("Couldn't load symbol for 'vkResetDescriptorPool': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    descriptor_pool,
    flags)
}


type VkAllocateDescriptorSets = fn (     C.Device,     &DescriptorSetAllocateInfo,     &C.DescriptorSet) Result

pub fn allocate_descriptor_sets(
    device                                          C.Device,
    p_allocate_info                                 &DescriptorSetAllocateInfo,
    p_descriptor_sets                               &C.DescriptorSet) Result {
      f := VkAllocateDescriptorSets((*loader_p).get_sym('vkAllocateDescriptorSets'
    ) or { 
        println("Couldn't load symbol for 'vkAllocateDescriptorSets': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_allocate_info,
    p_descriptor_sets)
}


type VkFreeDescriptorSets = fn (     C.Device,     C.DescriptorPool,     u32,     &C.DescriptorSet) Result

pub fn free_descriptor_sets(
    device                                          C.Device,
    descriptor_pool                                 C.DescriptorPool,
    descriptor_set_count                            u32,
    p_descriptor_sets                               &C.DescriptorSet) Result {
      f := VkFreeDescriptorSets((*loader_p).get_sym('vkFreeDescriptorSets'
    ) or { 
        println("Couldn't load symbol for 'vkFreeDescriptorSets': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    descriptor_pool,
    descriptor_set_count,
    p_descriptor_sets)
}


type VkUpdateDescriptorSets = fn (     C.Device,     u32,     &WriteDescriptorSet,     u32,     &CopyDescriptorSet) 

pub fn update_descriptor_sets(
    device                                          C.Device,
    descriptor_write_count                          u32,
    p_descriptor_writes                             &WriteDescriptorSet,
    descriptor_copy_count                           u32,
    p_descriptor_copies                             &CopyDescriptorSet)  {
      f := VkUpdateDescriptorSets((*loader_p).get_sym('vkUpdateDescriptorSets'
    ) or { 
        println("Couldn't load symbol for 'vkUpdateDescriptorSets': ${err}")
        return 
    })
    f(
    device,
    descriptor_write_count,
    p_descriptor_writes,
    descriptor_copy_count,
    p_descriptor_copies)
}


type VkCreateFramebuffer = fn (     C.Device,     &FramebufferCreateInfo,     &AllocationCallbacks,     &C.Framebuffer) Result

pub fn create_framebuffer(
    device                                          C.Device,
    p_create_info                                   &FramebufferCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_framebuffer                                   &C.Framebuffer) Result {
      f := VkCreateFramebuffer((*loader_p).get_sym('vkCreateFramebuffer'
    ) or { 
        println("Couldn't load symbol for 'vkCreateFramebuffer': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_framebuffer)
}


type VkDestroyFramebuffer = fn (     C.Device,     C.Framebuffer,     &AllocationCallbacks) 

pub fn destroy_framebuffer(
    device                                          C.Device,
    framebuffer                                     C.Framebuffer,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyFramebuffer((*loader_p).get_sym('vkDestroyFramebuffer'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyFramebuffer': ${err}")
        return 
    })
    f(
    device,
    framebuffer,
    p_allocator)
}


type VkCreateRenderPass = fn (     C.Device,     &RenderPassCreateInfo,     &AllocationCallbacks,     &C.RenderPass) Result

pub fn create_render_pass(
    device                                          C.Device,
    p_create_info                                   &RenderPassCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_render_pass                                   &C.RenderPass) Result {
      f := VkCreateRenderPass((*loader_p).get_sym('vkCreateRenderPass'
    ) or { 
        println("Couldn't load symbol for 'vkCreateRenderPass': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_render_pass)
}


type VkDestroyRenderPass = fn (     C.Device,     C.RenderPass,     &AllocationCallbacks) 

pub fn destroy_render_pass(
    device                                          C.Device,
    render_pass                                     C.RenderPass,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyRenderPass((*loader_p).get_sym('vkDestroyRenderPass'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyRenderPass': ${err}")
        return 
    })
    f(
    device,
    render_pass,
    p_allocator)
}


type VkGetRenderAreaGranularity = fn (     C.Device,     C.RenderPass,     &Extent2D) 

pub fn get_render_area_granularity(
    device                                          C.Device,
    render_pass                                     C.RenderPass,
    p_granularity                                   &Extent2D)  {
      f := VkGetRenderAreaGranularity((*loader_p).get_sym('vkGetRenderAreaGranularity'
    ) or { 
        println("Couldn't load symbol for 'vkGetRenderAreaGranularity': ${err}")
        return 
    })
    f(
    device,
    render_pass,
    p_granularity)
}


type VkCreateCommandPool = fn (     C.Device,     &CommandPoolCreateInfo,     &AllocationCallbacks,     &C.CommandPool) Result

pub fn create_command_pool(
    device                                          C.Device,
    p_create_info                                   &CommandPoolCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_command_pool                                  &C.CommandPool) Result {
      f := VkCreateCommandPool((*loader_p).get_sym('vkCreateCommandPool'
    ) or { 
        println("Couldn't load symbol for 'vkCreateCommandPool': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_command_pool)
}


type VkDestroyCommandPool = fn (     C.Device,     C.CommandPool,     &AllocationCallbacks) 

pub fn destroy_command_pool(
    device                                          C.Device,
    command_pool                                    C.CommandPool,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyCommandPool((*loader_p).get_sym('vkDestroyCommandPool'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyCommandPool': ${err}")
        return 
    })
    f(
    device,
    command_pool,
    p_allocator)
}


type VkResetCommandPool = fn (     C.Device,     C.CommandPool,     CommandPoolResetFlags) Result

pub fn reset_command_pool(
    device                                          C.Device,
    command_pool                                    C.CommandPool,
    flags                                           CommandPoolResetFlags) Result {
      f := VkResetCommandPool((*loader_p).get_sym('vkResetCommandPool'
    ) or { 
        println("Couldn't load symbol for 'vkResetCommandPool': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    command_pool,
    flags)
}


type VkAllocateCommandBuffers = fn (     C.Device,     &CommandBufferAllocateInfo,     &C.CommandBuffer) Result

pub fn allocate_command_buffers(
    device                                          C.Device,
    p_allocate_info                                 &CommandBufferAllocateInfo,
    p_command_buffers                               &C.CommandBuffer) Result {
      f := VkAllocateCommandBuffers((*loader_p).get_sym('vkAllocateCommandBuffers'
    ) or { 
        println("Couldn't load symbol for 'vkAllocateCommandBuffers': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_allocate_info,
    p_command_buffers)
}


type VkFreeCommandBuffers = fn (     C.Device,     C.CommandPool,     u32,     &C.CommandBuffer) 

pub fn free_command_buffers(
    device                                          C.Device,
    command_pool                                    C.CommandPool,
    command_buffer_count                            u32,
    p_command_buffers                               &C.CommandBuffer)  {
      f := VkFreeCommandBuffers((*loader_p).get_sym('vkFreeCommandBuffers'
    ) or { 
        println("Couldn't load symbol for 'vkFreeCommandBuffers': ${err}")
        return 
    })
    f(
    device,
    command_pool,
    command_buffer_count,
    p_command_buffers)
}


type VkBeginCommandBuffer = fn (     C.CommandBuffer,     &CommandBufferBeginInfo) Result

pub fn begin_command_buffer(
    command_buffer                                  C.CommandBuffer,
    p_begin_info                                    &CommandBufferBeginInfo) Result {
      f := VkBeginCommandBuffer((*loader_p).get_sym('vkBeginCommandBuffer'
    ) or { 
        println("Couldn't load symbol for 'vkBeginCommandBuffer': ${err}")
        return Result.error_unknown
    })
    return f(
    command_buffer,
    p_begin_info)
}


type VkEndCommandBuffer = fn (     C.CommandBuffer) Result

pub fn end_command_buffer(
    command_buffer                                  C.CommandBuffer) Result {
      f := VkEndCommandBuffer((*loader_p).get_sym('vkEndCommandBuffer'
    ) or { 
        println("Couldn't load symbol for 'vkEndCommandBuffer': ${err}")
        return Result.error_unknown
    })
    return f(
    command_buffer)
}


type VkResetCommandBuffer = fn (     C.CommandBuffer,     CommandBufferResetFlags) Result

pub fn reset_command_buffer(
    command_buffer                                  C.CommandBuffer,
    flags                                           CommandBufferResetFlags) Result {
      f := VkResetCommandBuffer((*loader_p).get_sym('vkResetCommandBuffer'
    ) or { 
        println("Couldn't load symbol for 'vkResetCommandBuffer': ${err}")
        return Result.error_unknown
    })
    return f(
    command_buffer,
    flags)
}


type VkCmdBindPipeline = fn (     C.CommandBuffer,     PipelineBindPoint,     C.Pipeline) 

pub fn cmd_bind_pipeline(
    command_buffer                                  C.CommandBuffer,
    pipeline_bind_point                             PipelineBindPoint,
    pipeline                                        C.Pipeline)  {
      f := VkCmdBindPipeline((*loader_p).get_sym('vkCmdBindPipeline'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindPipeline': ${err}")
        return 
    })
    f(
    command_buffer,
    pipeline_bind_point,
    pipeline)
}


type VkCmdSetViewport = fn (     C.CommandBuffer,     u32,     u32,     &Viewport) 

pub fn cmd_set_viewport(
    command_buffer                                  C.CommandBuffer,
    first_viewport                                  u32,
    viewport_count                                  u32,
    p_viewports                                     &Viewport)  {
      f := VkCmdSetViewport((*loader_p).get_sym('vkCmdSetViewport'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetViewport': ${err}")
        return 
    })
    f(
    command_buffer,
    first_viewport,
    viewport_count,
    p_viewports)
}


type VkCmdSetScissor = fn (     C.CommandBuffer,     u32,     u32,     &Rect2D) 

pub fn cmd_set_scissor(
    command_buffer                                  C.CommandBuffer,
    first_scissor                                   u32,
    scissor_count                                   u32,
    p_scissors                                      &Rect2D)  {
      f := VkCmdSetScissor((*loader_p).get_sym('vkCmdSetScissor'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetScissor': ${err}")
        return 
    })
    f(
    command_buffer,
    first_scissor,
    scissor_count,
    p_scissors)
}


type VkCmdSetLineWidth = fn (     C.CommandBuffer,     f32) 

pub fn cmd_set_line_width(
    command_buffer                                  C.CommandBuffer,
    line_width                                      f32)  {
      f := VkCmdSetLineWidth((*loader_p).get_sym('vkCmdSetLineWidth'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetLineWidth': ${err}")
        return 
    })
    f(
    command_buffer,
    line_width)
}


type VkCmdSetDepthBias = fn (     C.CommandBuffer,     f32,     f32,     f32) 

pub fn cmd_set_depth_bias(
    command_buffer                                  C.CommandBuffer,
    depth_bias_constant_factor                      f32,
    depth_bias_clamp                                f32,
    depth_bias_slope_factor                         f32)  {
      f := VkCmdSetDepthBias((*loader_p).get_sym('vkCmdSetDepthBias'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthBias': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_bias_constant_factor,
    depth_bias_clamp,
    depth_bias_slope_factor)
}


type VkCmdSetBlendConstants = fn (     C.CommandBuffer,     []f32) 

pub fn cmd_set_blend_constants(
    command_buffer                                  C.CommandBuffer,
    blend_constants                                 []f32)  {
      f := VkCmdSetBlendConstants((*loader_p).get_sym('vkCmdSetBlendConstants'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetBlendConstants': ${err}")
        return 
    })
    f(
    command_buffer,
    blend_constants)
}


type VkCmdSetDepthBounds = fn (     C.CommandBuffer,     f32,     f32) 

pub fn cmd_set_depth_bounds(
    command_buffer                                  C.CommandBuffer,
    min_depth_bounds                                f32,
    max_depth_bounds                                f32)  {
      f := VkCmdSetDepthBounds((*loader_p).get_sym('vkCmdSetDepthBounds'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthBounds': ${err}")
        return 
    })
    f(
    command_buffer,
    min_depth_bounds,
    max_depth_bounds)
}


type VkCmdSetStencilCompareMask = fn (     C.CommandBuffer,     StencilFaceFlags,     u32) 

pub fn cmd_set_stencil_compare_mask(
    command_buffer                                  C.CommandBuffer,
    face_mask                                       StencilFaceFlags,
    compare_mask                                    u32)  {
      f := VkCmdSetStencilCompareMask((*loader_p).get_sym('vkCmdSetStencilCompareMask'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetStencilCompareMask': ${err}")
        return 
    })
    f(
    command_buffer,
    face_mask,
    compare_mask)
}


type VkCmdSetStencilWriteMask = fn (     C.CommandBuffer,     StencilFaceFlags,     u32) 

pub fn cmd_set_stencil_write_mask(
    command_buffer                                  C.CommandBuffer,
    face_mask                                       StencilFaceFlags,
    write_mask                                      u32)  {
      f := VkCmdSetStencilWriteMask((*loader_p).get_sym('vkCmdSetStencilWriteMask'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetStencilWriteMask': ${err}")
        return 
    })
    f(
    command_buffer,
    face_mask,
    write_mask)
}


type VkCmdSetStencilReference = fn (     C.CommandBuffer,     StencilFaceFlags,     u32) 

pub fn cmd_set_stencil_reference(
    command_buffer                                  C.CommandBuffer,
    face_mask                                       StencilFaceFlags,
    reference                                       u32)  {
      f := VkCmdSetStencilReference((*loader_p).get_sym('vkCmdSetStencilReference'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetStencilReference': ${err}")
        return 
    })
    f(
    command_buffer,
    face_mask,
    reference)
}


type VkCmdBindDescriptorSets = fn (     C.CommandBuffer,     PipelineBindPoint,     C.PipelineLayout,     u32,     u32,     &C.DescriptorSet,     u32,     &u32) 

pub fn cmd_bind_descriptor_sets(
    command_buffer                                  C.CommandBuffer,
    pipeline_bind_point                             PipelineBindPoint,
    layout                                          C.PipelineLayout,
    first_set                                       u32,
    descriptor_set_count                            u32,
    p_descriptor_sets                               &C.DescriptorSet,
    dynamic_offset_count                            u32,
    p_dynamic_offsets                               &u32)  {
      f := VkCmdBindDescriptorSets((*loader_p).get_sym('vkCmdBindDescriptorSets'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindDescriptorSets': ${err}")
        return 
    })
    f(
    command_buffer,
    pipeline_bind_point,
    layout,
    first_set,
    descriptor_set_count,
    p_descriptor_sets,
    dynamic_offset_count,
    p_dynamic_offsets)
}


type VkCmdBindIndexBuffer = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     IndexType) 

pub fn cmd_bind_index_buffer(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    index_type                                      IndexType)  {
      f := VkCmdBindIndexBuffer((*loader_p).get_sym('vkCmdBindIndexBuffer'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindIndexBuffer': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    index_type)
}


type VkCmdBindVertexBuffers = fn (     C.CommandBuffer,     u32,     u32,     &C.Buffer,     &DeviceSize) 

pub fn cmd_bind_vertex_buffers(
    command_buffer                                  C.CommandBuffer,
    first_binding                                   u32,
    binding_count                                   u32,
    p_buffers                                       &C.Buffer,
    p_offsets                                       &DeviceSize)  {
      f := VkCmdBindVertexBuffers((*loader_p).get_sym('vkCmdBindVertexBuffers'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindVertexBuffers': ${err}")
        return 
    })
    f(
    command_buffer,
    first_binding,
    binding_count,
    p_buffers,
    p_offsets)
}


type VkCmdDraw = fn (     C.CommandBuffer,     u32,     u32,     u32,     u32) 

pub fn cmd_draw(
    command_buffer                                  C.CommandBuffer,
    vertex_count                                    u32,
    instance_count                                  u32,
    first_vertex                                    u32,
    first_instance                                  u32)  {
      f := VkCmdDraw((*loader_p).get_sym('vkCmdDraw'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDraw': ${err}")
        return 
    })
    f(
    command_buffer,
    vertex_count,
    instance_count,
    first_vertex,
    first_instance)
}


type VkCmdDrawIndexed = fn (     C.CommandBuffer,     u32,     u32,     u32,     i32,     u32) 

pub fn cmd_draw_indexed(
    command_buffer                                  C.CommandBuffer,
    index_count                                     u32,
    instance_count                                  u32,
    first_index                                     u32,
    vertex_offset                                   i32,
    first_instance                                  u32)  {
      f := VkCmdDrawIndexed((*loader_p).get_sym('vkCmdDrawIndexed'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawIndexed': ${err}")
        return 
    })
    f(
    command_buffer,
    index_count,
    instance_count,
    first_index,
    vertex_offset,
    first_instance)
}


type VkCmdDrawIndirect = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_indirect(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    draw_count                                      u32,
    stride                                          u32)  {
      f := VkCmdDrawIndirect((*loader_p).get_sym('vkCmdDrawIndirect'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawIndirect': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    draw_count,
    stride)
}


type VkCmdDrawIndexedIndirect = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_indexed_indirect(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    draw_count                                      u32,
    stride                                          u32)  {
      f := VkCmdDrawIndexedIndirect((*loader_p).get_sym('vkCmdDrawIndexedIndirect'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawIndexedIndirect': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    draw_count,
    stride)
}


type VkCmdDispatch = fn (     C.CommandBuffer,     u32,     u32,     u32) 

pub fn cmd_dispatch(
    command_buffer                                  C.CommandBuffer,
    group_count_x                                   u32,
    group_count_y                                   u32,
    group_count_z                                   u32)  {
      f := VkCmdDispatch((*loader_p).get_sym('vkCmdDispatch'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDispatch': ${err}")
        return 
    })
    f(
    command_buffer,
    group_count_x,
    group_count_y,
    group_count_z)
}


type VkCmdDispatchIndirect = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize) 

pub fn cmd_dispatch_indirect(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize)  {
      f := VkCmdDispatchIndirect((*loader_p).get_sym('vkCmdDispatchIndirect'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDispatchIndirect': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset)
}


type VkCmdCopyBuffer = fn (     C.CommandBuffer,     C.Buffer,     C.Buffer,     u32,     &BufferCopy) 

pub fn cmd_copy_buffer(
    command_buffer                                  C.CommandBuffer,
    src_buffer                                      C.Buffer,
    dst_buffer                                      C.Buffer,
    region_count                                    u32,
    p_regions                                       &BufferCopy)  {
      f := VkCmdCopyBuffer((*loader_p).get_sym('vkCmdCopyBuffer'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyBuffer': ${err}")
        return 
    })
    f(
    command_buffer,
    src_buffer,
    dst_buffer,
    region_count,
    p_regions)
}


type VkCmdCopyImage = fn (     C.CommandBuffer,     C.Image,     ImageLayout,     C.Image,     ImageLayout,     u32,     &ImageCopy) 

pub fn cmd_copy_image(
    command_buffer                                  C.CommandBuffer,
    src_image                                       C.Image,
    src_image_layout                                ImageLayout,
    dst_image                                       C.Image,
    dst_image_layout                                ImageLayout,
    region_count                                    u32,
    p_regions                                       &ImageCopy)  {
      f := VkCmdCopyImage((*loader_p).get_sym('vkCmdCopyImage'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyImage': ${err}")
        return 
    })
    f(
    command_buffer,
    src_image,
    src_image_layout,
    dst_image,
    dst_image_layout,
    region_count,
    p_regions)
}


type VkCmdBlitImage = fn (     C.CommandBuffer,     C.Image,     ImageLayout,     C.Image,     ImageLayout,     u32,     &ImageBlit,     Filter) 

pub fn cmd_blit_image(
    command_buffer                                  C.CommandBuffer,
    src_image                                       C.Image,
    src_image_layout                                ImageLayout,
    dst_image                                       C.Image,
    dst_image_layout                                ImageLayout,
    region_count                                    u32,
    p_regions                                       &ImageBlit,
    filter                                          Filter)  {
      f := VkCmdBlitImage((*loader_p).get_sym('vkCmdBlitImage'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBlitImage': ${err}")
        return 
    })
    f(
    command_buffer,
    src_image,
    src_image_layout,
    dst_image,
    dst_image_layout,
    region_count,
    p_regions,
    filter)
}


type VkCmdCopyBufferToImage = fn (     C.CommandBuffer,     C.Buffer,     C.Image,     ImageLayout,     u32,     &BufferImageCopy) 

pub fn cmd_copy_buffer_to_image(
    command_buffer                                  C.CommandBuffer,
    src_buffer                                      C.Buffer,
    dst_image                                       C.Image,
    dst_image_layout                                ImageLayout,
    region_count                                    u32,
    p_regions                                       &BufferImageCopy)  {
      f := VkCmdCopyBufferToImage((*loader_p).get_sym('vkCmdCopyBufferToImage'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyBufferToImage': ${err}")
        return 
    })
    f(
    command_buffer,
    src_buffer,
    dst_image,
    dst_image_layout,
    region_count,
    p_regions)
}


type VkCmdCopyImageToBuffer = fn (     C.CommandBuffer,     C.Image,     ImageLayout,     C.Buffer,     u32,     &BufferImageCopy) 

pub fn cmd_copy_image_to_buffer(
    command_buffer                                  C.CommandBuffer,
    src_image                                       C.Image,
    src_image_layout                                ImageLayout,
    dst_buffer                                      C.Buffer,
    region_count                                    u32,
    p_regions                                       &BufferImageCopy)  {
      f := VkCmdCopyImageToBuffer((*loader_p).get_sym('vkCmdCopyImageToBuffer'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyImageToBuffer': ${err}")
        return 
    })
    f(
    command_buffer,
    src_image,
    src_image_layout,
    dst_buffer,
    region_count,
    p_regions)
}


type VkCmdUpdateBuffer = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     DeviceSize,     voidptr) 

pub fn cmd_update_buffer(
    command_buffer                                  C.CommandBuffer,
    dst_buffer                                      C.Buffer,
    dst_offset                                      DeviceSize,
    data_size                                       DeviceSize,
    p_data                                          voidptr)  {
      f := VkCmdUpdateBuffer((*loader_p).get_sym('vkCmdUpdateBuffer'
    ) or { 
        println("Couldn't load symbol for 'vkCmdUpdateBuffer': ${err}")
        return 
    })
    f(
    command_buffer,
    dst_buffer,
    dst_offset,
    data_size,
    p_data)
}


type VkCmdFillBuffer = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     DeviceSize,     u32) 

pub fn cmd_fill_buffer(
    command_buffer                                  C.CommandBuffer,
    dst_buffer                                      C.Buffer,
    dst_offset                                      DeviceSize,
    size                                            DeviceSize,
    data                                            u32)  {
      f := VkCmdFillBuffer((*loader_p).get_sym('vkCmdFillBuffer'
    ) or { 
        println("Couldn't load symbol for 'vkCmdFillBuffer': ${err}")
        return 
    })
    f(
    command_buffer,
    dst_buffer,
    dst_offset,
    size,
    data)
}


type VkCmdClearColorImage = fn (     C.CommandBuffer,     C.Image,     ImageLayout,     &ClearColorValue,     u32,     &ImageSubresourceRange) 

pub fn cmd_clear_color_image(
    command_buffer                                  C.CommandBuffer,
    image                                           C.Image,
    image_layout                                    ImageLayout,
    p_color                                         &ClearColorValue,
    range_count                                     u32,
    p_ranges                                        &ImageSubresourceRange)  {
      f := VkCmdClearColorImage((*loader_p).get_sym('vkCmdClearColorImage'
    ) or { 
        println("Couldn't load symbol for 'vkCmdClearColorImage': ${err}")
        return 
    })
    f(
    command_buffer,
    image,
    image_layout,
    p_color,
    range_count,
    p_ranges)
}


type VkCmdClearDepthStencilImage = fn (     C.CommandBuffer,     C.Image,     ImageLayout,     &ClearDepthStencilValue,     u32,     &ImageSubresourceRange) 

pub fn cmd_clear_depth_stencil_image(
    command_buffer                                  C.CommandBuffer,
    image                                           C.Image,
    image_layout                                    ImageLayout,
    p_depth_stencil                                 &ClearDepthStencilValue,
    range_count                                     u32,
    p_ranges                                        &ImageSubresourceRange)  {
      f := VkCmdClearDepthStencilImage((*loader_p).get_sym('vkCmdClearDepthStencilImage'
    ) or { 
        println("Couldn't load symbol for 'vkCmdClearDepthStencilImage': ${err}")
        return 
    })
    f(
    command_buffer,
    image,
    image_layout,
    p_depth_stencil,
    range_count,
    p_ranges)
}


type VkCmdClearAttachments = fn (     C.CommandBuffer,     u32,     &ClearAttachment,     u32,     &ClearRect) 

pub fn cmd_clear_attachments(
    command_buffer                                  C.CommandBuffer,
    attachment_count                                u32,
    p_attachments                                   &ClearAttachment,
    rect_count                                      u32,
    p_rects                                         &ClearRect)  {
      f := VkCmdClearAttachments((*loader_p).get_sym('vkCmdClearAttachments'
    ) or { 
        println("Couldn't load symbol for 'vkCmdClearAttachments': ${err}")
        return 
    })
    f(
    command_buffer,
    attachment_count,
    p_attachments,
    rect_count,
    p_rects)
}


type VkCmdResolveImage = fn (     C.CommandBuffer,     C.Image,     ImageLayout,     C.Image,     ImageLayout,     u32,     &ImageResolve) 

pub fn cmd_resolve_image(
    command_buffer                                  C.CommandBuffer,
    src_image                                       C.Image,
    src_image_layout                                ImageLayout,
    dst_image                                       C.Image,
    dst_image_layout                                ImageLayout,
    region_count                                    u32,
    p_regions                                       &ImageResolve)  {
      f := VkCmdResolveImage((*loader_p).get_sym('vkCmdResolveImage'
    ) or { 
        println("Couldn't load symbol for 'vkCmdResolveImage': ${err}")
        return 
    })
    f(
    command_buffer,
    src_image,
    src_image_layout,
    dst_image,
    dst_image_layout,
    region_count,
    p_regions)
}


type VkCmdSetEvent = fn (     C.CommandBuffer,     C.Event,     PipelineStageFlags) 

pub fn cmd_set_event(
    command_buffer                                  C.CommandBuffer,
    event                                           C.Event,
    stage_mask                                      PipelineStageFlags)  {
      f := VkCmdSetEvent((*loader_p).get_sym('vkCmdSetEvent'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetEvent': ${err}")
        return 
    })
    f(
    command_buffer,
    event,
    stage_mask)
}


type VkCmdResetEvent = fn (     C.CommandBuffer,     C.Event,     PipelineStageFlags) 

pub fn cmd_reset_event(
    command_buffer                                  C.CommandBuffer,
    event                                           C.Event,
    stage_mask                                      PipelineStageFlags)  {
      f := VkCmdResetEvent((*loader_p).get_sym('vkCmdResetEvent'
    ) or { 
        println("Couldn't load symbol for 'vkCmdResetEvent': ${err}")
        return 
    })
    f(
    command_buffer,
    event,
    stage_mask)
}


type VkCmdWaitEvents = fn (     C.CommandBuffer,     u32,     &C.Event,     PipelineStageFlags,     PipelineStageFlags,     u32,     &MemoryBarrier,     u32,     &BufferMemoryBarrier,     u32,     &ImageMemoryBarrier) 

pub fn cmd_wait_events(
    command_buffer                                  C.CommandBuffer,
    event_count                                     u32,
    p_events                                        &C.Event,
    src_stage_mask                                  PipelineStageFlags,
    dst_stage_mask                                  PipelineStageFlags,
    memory_barrier_count                            u32,
    p_memory_barriers                               &MemoryBarrier,
    buffer_memory_barrier_count                     u32,
    p_buffer_memory_barriers                        &BufferMemoryBarrier,
    image_memory_barrier_count                      u32,
    p_image_memory_barriers                         &ImageMemoryBarrier)  {
      f := VkCmdWaitEvents((*loader_p).get_sym('vkCmdWaitEvents'
    ) or { 
        println("Couldn't load symbol for 'vkCmdWaitEvents': ${err}")
        return 
    })
    f(
    command_buffer,
    event_count,
    p_events,
    src_stage_mask,
    dst_stage_mask,
    memory_barrier_count,
    p_memory_barriers,
    buffer_memory_barrier_count,
    p_buffer_memory_barriers,
    image_memory_barrier_count,
    p_image_memory_barriers)
}


type VkCmdPipelineBarrier = fn (     C.CommandBuffer,     PipelineStageFlags,     PipelineStageFlags,     DependencyFlags,     u32,     &MemoryBarrier,     u32,     &BufferMemoryBarrier,     u32,     &ImageMemoryBarrier) 

pub fn cmd_pipeline_barrier(
    command_buffer                                  C.CommandBuffer,
    src_stage_mask                                  PipelineStageFlags,
    dst_stage_mask                                  PipelineStageFlags,
    dependency_flags                                DependencyFlags,
    memory_barrier_count                            u32,
    p_memory_barriers                               &MemoryBarrier,
    buffer_memory_barrier_count                     u32,
    p_buffer_memory_barriers                        &BufferMemoryBarrier,
    image_memory_barrier_count                      u32,
    p_image_memory_barriers                         &ImageMemoryBarrier)  {
      f := VkCmdPipelineBarrier((*loader_p).get_sym('vkCmdPipelineBarrier'
    ) or { 
        println("Couldn't load symbol for 'vkCmdPipelineBarrier': ${err}")
        return 
    })
    f(
    command_buffer,
    src_stage_mask,
    dst_stage_mask,
    dependency_flags,
    memory_barrier_count,
    p_memory_barriers,
    buffer_memory_barrier_count,
    p_buffer_memory_barriers,
    image_memory_barrier_count,
    p_image_memory_barriers)
}


type VkCmdBeginQuery = fn (     C.CommandBuffer,     C.QueryPool,     u32,     QueryControlFlags) 

pub fn cmd_begin_query(
    command_buffer                                  C.CommandBuffer,
    query_pool                                      C.QueryPool,
    query                                           u32,
    flags                                           QueryControlFlags)  {
      f := VkCmdBeginQuery((*loader_p).get_sym('vkCmdBeginQuery'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBeginQuery': ${err}")
        return 
    })
    f(
    command_buffer,
    query_pool,
    query,
    flags)
}


type VkCmdEndQuery = fn (     C.CommandBuffer,     C.QueryPool,     u32) 

pub fn cmd_end_query(
    command_buffer                                  C.CommandBuffer,
    query_pool                                      C.QueryPool,
    query                                           u32)  {
      f := VkCmdEndQuery((*loader_p).get_sym('vkCmdEndQuery'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEndQuery': ${err}")
        return 
    })
    f(
    command_buffer,
    query_pool,
    query)
}


type VkCmdResetQueryPool = fn (     C.CommandBuffer,     C.QueryPool,     u32,     u32) 

pub fn cmd_reset_query_pool(
    command_buffer                                  C.CommandBuffer,
    query_pool                                      C.QueryPool,
    first_query                                     u32,
    query_count                                     u32)  {
      f := VkCmdResetQueryPool((*loader_p).get_sym('vkCmdResetQueryPool'
    ) or { 
        println("Couldn't load symbol for 'vkCmdResetQueryPool': ${err}")
        return 
    })
    f(
    command_buffer,
    query_pool,
    first_query,
    query_count)
}


type VkCmdWriteTimestamp = fn (     C.CommandBuffer,     PipelineStageFlagBits,     C.QueryPool,     u32) 

pub fn cmd_write_timestamp(
    command_buffer                                  C.CommandBuffer,
    pipeline_stage                                  PipelineStageFlagBits,
    query_pool                                      C.QueryPool,
    query                                           u32)  {
      f := VkCmdWriteTimestamp((*loader_p).get_sym('vkCmdWriteTimestamp'
    ) or { 
        println("Couldn't load symbol for 'vkCmdWriteTimestamp': ${err}")
        return 
    })
    f(
    command_buffer,
    pipeline_stage,
    query_pool,
    query)
}


type VkCmdCopyQueryPoolResults = fn (     C.CommandBuffer,     C.QueryPool,     u32,     u32,     C.Buffer,     DeviceSize,     DeviceSize,     QueryResultFlags) 

pub fn cmd_copy_query_pool_results(
    command_buffer                                  C.CommandBuffer,
    query_pool                                      C.QueryPool,
    first_query                                     u32,
    query_count                                     u32,
    dst_buffer                                      C.Buffer,
    dst_offset                                      DeviceSize,
    stride                                          DeviceSize,
    flags                                           QueryResultFlags)  {
      f := VkCmdCopyQueryPoolResults((*loader_p).get_sym('vkCmdCopyQueryPoolResults'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyQueryPoolResults': ${err}")
        return 
    })
    f(
    command_buffer,
    query_pool,
    first_query,
    query_count,
    dst_buffer,
    dst_offset,
    stride,
    flags)
}


type VkCmdPushConstants = fn (     C.CommandBuffer,     C.PipelineLayout,     ShaderStageFlags,     u32,     u32,     voidptr) 

pub fn cmd_push_constants(
    command_buffer                                  C.CommandBuffer,
    layout                                          C.PipelineLayout,
    stage_flags                                     ShaderStageFlags,
    offset                                          u32,
    size                                            u32,
    p_values                                        voidptr)  {
      f := VkCmdPushConstants((*loader_p).get_sym('vkCmdPushConstants'
    ) or { 
        println("Couldn't load symbol for 'vkCmdPushConstants': ${err}")
        return 
    })
    f(
    command_buffer,
    layout,
    stage_flags,
    offset,
    size,
    p_values)
}


type VkCmdBeginRenderPass = fn (     C.CommandBuffer,     &RenderPassBeginInfo,     SubpassContents) 

pub fn cmd_begin_render_pass(
    command_buffer                                  C.CommandBuffer,
    p_render_pass_begin                             &RenderPassBeginInfo,
    contents                                        SubpassContents)  {
      f := VkCmdBeginRenderPass((*loader_p).get_sym('vkCmdBeginRenderPass'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBeginRenderPass': ${err}")
        return 
    })
    f(
    command_buffer,
    p_render_pass_begin,
    contents)
}


type VkCmdNextSubpass = fn (     C.CommandBuffer,     SubpassContents) 

pub fn cmd_next_subpass(
    command_buffer                                  C.CommandBuffer,
    contents                                        SubpassContents)  {
      f := VkCmdNextSubpass((*loader_p).get_sym('vkCmdNextSubpass'
    ) or { 
        println("Couldn't load symbol for 'vkCmdNextSubpass': ${err}")
        return 
    })
    f(
    command_buffer,
    contents)
}


type VkCmdEndRenderPass = fn (     C.CommandBuffer) 

pub fn cmd_end_render_pass(
    command_buffer                                  C.CommandBuffer)  {
      f := VkCmdEndRenderPass((*loader_p).get_sym('vkCmdEndRenderPass'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEndRenderPass': ${err}")
        return 
    })
    f(
    command_buffer)
}


type VkCmdExecuteCommands = fn (     C.CommandBuffer,     u32,     &C.CommandBuffer) 

pub fn cmd_execute_commands(
    command_buffer                                  C.CommandBuffer,
    command_buffer_count                            u32,
    p_command_buffers                               &C.CommandBuffer)  {
      f := VkCmdExecuteCommands((*loader_p).get_sym('vkCmdExecuteCommands'
    ) or { 
        println("Couldn't load symbol for 'vkCmdExecuteCommands': ${err}")
        return 
    })
    f(
    command_buffer,
    command_buffer_count,
    p_command_buffers)
}




// VK_VERSION_1_1 is a preprocessor guard. Do not pass it to API calls.
const version_1_1 = 1
// Vulkan 1.1 version number
pub const api_version_1_1 = make_api_version(0, 1, 1, 0)// Patch version should always be set to 0

pub type C.SamplerYcbcrConversion = voidptr
pub type C.DescriptorUpdateTemplate = voidptr
pub const max_device_group_size             = u32(32)
pub const luid_size                         = u32(8)
pub const queue_family_external             = ~u32(1)

pub enum PointClippingBehavior {
    point_clipping_behavior_all_clip_planes = int(0)
    point_clipping_behavior_user_clip_planes_only = int(1)
    point_clipping_behavior_max_enum = int(0x7FFFFFFF)
}


pub enum TessellationDomainOrigin {
    tessellation_domain_origin_upper_left = int(0)
    tessellation_domain_origin_lower_left = int(1)
    tessellation_domain_origin_max_enum = int(0x7FFFFFFF)
}


pub enum SamplerYcbcrModelConversion {
    sampler_ycbcr_model_conversion_rgb_identity = int(0)
    sampler_ycbcr_model_conversion_ycbcr_identity = int(1)
    sampler_ycbcr_model_conversion_ycbcr_709 = int(2)
    sampler_ycbcr_model_conversion_ycbcr_601 = int(3)
    sampler_ycbcr_model_conversion_ycbcr_2020 = int(4)
    sampler_ycbcr_model_conversion_max_enum = int(0x7FFFFFFF)
}


pub enum SamplerYcbcrRange {
    sampler_ycbcr_range_itu_full = int(0)
    sampler_ycbcr_range_itu_narrow = int(1)
    sampler_ycbcr_range_max_enum = int(0x7FFFFFFF)
}


pub enum ChromaLocation {
    chroma_location_cosited_even = int(0)
    chroma_location_midpoint = int(1)
    chroma_location_max_enum = int(0x7FFFFFFF)
}


pub enum DescriptorUpdateTemplateType {
    descriptor_update_template_type_descriptor_set = int(0)
    descriptor_update_template_type_push_descriptors_khr = int(1)
    descriptor_update_template_type_max_enum = int(0x7FFFFFFF)
}


pub enum SubgroupFeatureFlagBits {
    subgroup_feature_basic_bit = int(0x00000001)
    subgroup_feature_vote_bit = int(0x00000002)
    subgroup_feature_arithmetic_bit = int(0x00000004)
    subgroup_feature_ballot_bit = int(0x00000008)
    subgroup_feature_shuffle_bit = int(0x00000010)
    subgroup_feature_shuffle_relative_bit = int(0x00000020)
    subgroup_feature_clustered_bit = int(0x00000040)
    subgroup_feature_quad_bit = int(0x00000080)
    subgroup_feature_partitioned_bit_nv = int(0x00000100)
    subgroup_feature_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type SubgroupFeatureFlags = u32

pub enum PeerMemoryFeatureFlagBits {
    peer_memory_feature_copy_src_bit = int(0x00000001)
    peer_memory_feature_copy_dst_bit = int(0x00000002)
    peer_memory_feature_generic_src_bit = int(0x00000004)
    peer_memory_feature_generic_dst_bit = int(0x00000008)
    peer_memory_feature_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type PeerMemoryFeatureFlags = u32

pub enum MemoryAllocateFlagBits {
    memory_allocate_device_mask_bit = int(0x00000001)
    memory_allocate_device_address_bit = int(0x00000002)
    memory_allocate_device_address_capture_replay_bit = int(0x00000004)
    memory_allocate_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type MemoryAllocateFlags = u32
pub type CommandPoolTrimFlags = u32
pub type DescriptorUpdateTemplateCreateFlags = u32

pub enum ExternalMemoryHandleTypeFlagBits {
    external_memory_handle_type_opaque_fd_bit = int(0x00000001)
    external_memory_handle_type_opaque_win32_bit = int(0x00000002)
    external_memory_handle_type_opaque_win32_kmt_bit = int(0x00000004)
    external_memory_handle_type_d3d11_texture_bit = int(0x00000008)
    external_memory_handle_type_d3d11_texture_kmt_bit = int(0x00000010)
    external_memory_handle_type_d3d12_heap_bit = int(0x00000020)
    external_memory_handle_type_d3d12_resource_bit = int(0x00000040)
    external_memory_handle_type_dma_buf_bit_ext = int(0x00000200)
    external_memory_handle_type_android_hardware_buffer_bit_android = int(0x00000400)
    external_memory_handle_type_host_allocation_bit_ext = int(0x00000080)
    external_memory_handle_type_host_mapped_foreign_memory_bit_ext = int(0x00000100)
    external_memory_handle_type_zircon_vmo_bit_fuchsia = int(0x00000800)
    external_memory_handle_type_rdma_address_bit_nv = int(0x00001000)
    external_memory_handle_type_screen_buffer_bit_qnx = int(0x00004000)
    external_memory_handle_type_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ExternalMemoryHandleTypeFlags = u32

pub enum ExternalMemoryFeatureFlagBits {
    external_memory_feature_dedicated_only_bit = int(0x00000001)
    external_memory_feature_exportable_bit = int(0x00000002)
    external_memory_feature_importable_bit = int(0x00000004)
    external_memory_feature_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ExternalMemoryFeatureFlags = u32

pub enum ExternalFenceHandleTypeFlagBits {
    external_fence_handle_type_opaque_fd_bit = int(0x00000001)
    external_fence_handle_type_opaque_win32_bit = int(0x00000002)
    external_fence_handle_type_opaque_win32_kmt_bit = int(0x00000004)
    external_fence_handle_type_sync_fd_bit = int(0x00000008)
    external_fence_handle_type_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ExternalFenceHandleTypeFlags = u32

pub enum ExternalFenceFeatureFlagBits {
    external_fence_feature_exportable_bit = int(0x00000001)
    external_fence_feature_importable_bit = int(0x00000002)
    external_fence_feature_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ExternalFenceFeatureFlags = u32

pub enum FenceImportFlagBits {
    fence_import_temporary_bit = int(0x00000001)
    fence_import_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type FenceImportFlags = u32

pub enum SemaphoreImportFlagBits {
    semaphore_import_temporary_bit = int(0x00000001)
    semaphore_import_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type SemaphoreImportFlags = u32

pub enum ExternalSemaphoreHandleTypeFlagBits {
    external_semaphore_handle_type_opaque_fd_bit = int(0x00000001)
    external_semaphore_handle_type_opaque_win32_bit = int(0x00000002)
    external_semaphore_handle_type_opaque_win32_kmt_bit = int(0x00000004)
    external_semaphore_handle_type_d3d12_fence_bit = int(0x00000008)
    external_semaphore_handle_type_sync_fd_bit = int(0x00000010)
    external_semaphore_handle_type_zircon_event_bit_fuchsia = int(0x00000080)
    external_semaphore_handle_type_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ExternalSemaphoreHandleTypeFlags = u32

pub enum ExternalSemaphoreFeatureFlagBits {
    external_semaphore_feature_exportable_bit = int(0x00000001)
    external_semaphore_feature_importable_bit = int(0x00000002)
    external_semaphore_feature_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ExternalSemaphoreFeatureFlags = u32
// PhysicalDeviceSubgroupProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceSubgroupProperties {
mut:
    s_type                        StructureType
    p_next                        voidptr
    subgroup_size                 u32
    supported_stages              ShaderStageFlags
    supported_operations          SubgroupFeatureFlags
    quad_operations_in_all_stages Bool32
} 

pub struct BindBufferMemoryInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    buffer                 C.Buffer
    memory                 C.DeviceMemory
    memory_offset          DeviceSize
} 

pub struct BindImageMemoryInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image                  C.Image
    memory                 C.DeviceMemory
    memory_offset          DeviceSize
} 

// PhysicalDevice16BitStorageFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevice16BitStorageFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    storage_buffer16_bit_access Bool32
    uniform_and_storage_buffer16_bit_access Bool32
    storage_push_constant16 Bool32
    storage_input_output16 Bool32
} 

// MemoryDedicatedRequirements extends VkMemoryRequirements2
pub struct MemoryDedicatedRequirements {
mut:
    s_type                 StructureType
    p_next                 voidptr
    prefers_dedicated_allocation Bool32
    requires_dedicated_allocation Bool32
} 

// MemoryDedicatedAllocateInfo extends VkMemoryAllocateInfo
pub struct MemoryDedicatedAllocateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image                  C.Image
    buffer                 C.Buffer
} 

// MemoryAllocateFlagsInfo extends VkMemoryAllocateInfo
pub struct MemoryAllocateFlagsInfo {
mut:
    s_type                       StructureType
    p_next                       voidptr
    flags                        MemoryAllocateFlags
    device_mask                  u32
} 

// DeviceGroupRenderPassBeginInfo extends VkRenderPassBeginInfo,VkRenderingInfo
pub struct DeviceGroupRenderPassBeginInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_mask            u32
    device_render_area_count u32
    p_device_render_areas  &Rect2D
} 

// DeviceGroupCommandBufferBeginInfo extends VkCommandBufferBeginInfo
pub struct DeviceGroupCommandBufferBeginInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_mask            u32
} 

// DeviceGroupSubmitInfo extends VkSubmitInfo
pub struct DeviceGroupSubmitInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    wait_semaphore_count   u32
    p_wait_semaphore_device_indices &u32
    command_buffer_count   u32
    p_command_buffer_device_masks &u32
    signal_semaphore_count u32
    p_signal_semaphore_device_indices &u32
} 

// DeviceGroupBindSparseInfo extends VkBindSparseInfo
pub struct DeviceGroupBindSparseInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    resource_device_index  u32
    memory_device_index    u32
} 

// BindBufferMemoryDeviceGroupInfo extends VkBindBufferMemoryInfo
pub struct BindBufferMemoryDeviceGroupInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_index_count     u32
    p_device_indices       &u32
} 

// BindImageMemoryDeviceGroupInfo extends VkBindImageMemoryInfo
pub struct BindImageMemoryDeviceGroupInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_index_count     u32
    p_device_indices       &u32
    split_instance_bind_region_count u32
    p_split_instance_bind_regions &Rect2D
} 

pub struct PhysicalDeviceGroupProperties {
mut:
    s_type                  StructureType
    p_next                  voidptr
    physical_device_count   u32
    physical_devices        []C.PhysicalDevice
    subset_allocation       Bool32
} 

// DeviceGroupDeviceCreateInfo extends VkDeviceCreateInfo
pub struct DeviceGroupDeviceCreateInfo {
mut:
    s_type                         StructureType
    p_next                         voidptr
    physical_device_count          u32
    p_physical_devices             &C.PhysicalDevice
} 

pub struct BufferMemoryRequirementsInfo2 {
mut:
    s_type                 StructureType
    p_next                 voidptr
    buffer                 C.Buffer
} 

pub struct ImageMemoryRequirementsInfo2 {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image                  C.Image
} 

pub struct ImageSparseMemoryRequirementsInfo2 {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image                  C.Image
} 

pub struct MemoryRequirements2 {
mut:
    s_type                      StructureType
    p_next                      voidptr
    memory_requirements         MemoryRequirements
} 

pub struct SparseImageMemoryRequirements2 {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    memory_requirements                    SparseImageMemoryRequirements
} 

// PhysicalDeviceFeatures2 extends VkDeviceCreateInfo
pub struct PhysicalDeviceFeatures2 {
mut:
    s_type                          StructureType
    p_next                          voidptr
    features                        PhysicalDeviceFeatures
} 

pub struct PhysicalDeviceProperties2 {
mut:
    s_type                            StructureType
    p_next                            voidptr
    properties                        PhysicalDeviceProperties
} 

pub struct FormatProperties2 {
mut:
    s_type                    StructureType
    p_next                    voidptr
    format_properties         FormatProperties
} 

pub struct ImageFormatProperties2 {
mut:
    s_type                         StructureType
    p_next                         voidptr
    image_format_properties        ImageFormatProperties
} 

pub struct PhysicalDeviceImageFormatInfo2 {
mut:
    s_type                    StructureType
    p_next                    voidptr
    format                    Format
    vktype                    ImageType
    tiling                    ImageTiling
    usage                     ImageUsageFlags
    flags                     ImageCreateFlags
} 

pub struct QueueFamilyProperties2 {
mut:
    s_type                         StructureType
    p_next                         voidptr
    queue_family_properties        QueueFamilyProperties
} 

pub struct PhysicalDeviceMemoryProperties2 {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    memory_properties                       PhysicalDeviceMemoryProperties
} 

pub struct SparseImageFormatProperties2 {
mut:
    s_type                               StructureType
    p_next                               voidptr
    properties                           SparseImageFormatProperties
} 

pub struct PhysicalDeviceSparseImageFormatInfo2 {
mut:
    s_type                       StructureType
    p_next                       voidptr
    format                       Format
    vktype                       ImageType
    samples                      SampleCountFlagBits
    usage                        ImageUsageFlags
    tiling                       ImageTiling
} 

// PhysicalDevicePointClippingProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDevicePointClippingProperties {
mut:
    s_type                         StructureType
    p_next                         voidptr
    point_clipping_behavior        PointClippingBehavior
} 

pub struct InputAttachmentAspectReference {
mut:
    subpass                   u32
    input_attachment_index    u32
    aspect_mask               ImageAspectFlags
} 

// RenderPassInputAttachmentAspectCreateInfo extends VkRenderPassCreateInfo
pub struct RenderPassInputAttachmentAspectCreateInfo {
mut:
    s_type                                         StructureType
    p_next                                         voidptr
    aspect_reference_count                         u32
    p_aspect_references                            &InputAttachmentAspectReference
} 

// ImageViewUsageCreateInfo extends VkImageViewCreateInfo
pub struct ImageViewUsageCreateInfo {
mut:
    s_type                   StructureType
    p_next                   voidptr
    usage                    ImageUsageFlags
} 

// PipelineTessellationDomainOriginStateCreateInfo extends VkPipelineTessellationStateCreateInfo
pub struct PipelineTessellationDomainOriginStateCreateInfo {
mut:
    s_type                            StructureType
    p_next                            voidptr
    domain_origin                     TessellationDomainOrigin
} 

// RenderPassMultiviewCreateInfo extends VkRenderPassCreateInfo
pub struct RenderPassMultiviewCreateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    subpass_count          u32
    p_view_masks           &u32
    dependency_count       u32
    p_view_offsets         &i32
    correlation_mask_count u32
    p_correlation_masks    &u32
} 

// PhysicalDeviceMultiviewFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMultiviewFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    multiview              Bool32
    multiview_geometry_shader Bool32
    multiview_tessellation_shader Bool32
} 

// PhysicalDeviceMultiviewProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceMultiviewProperties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_multiview_view_count u32
    max_multiview_instance_index u32
} 

// PhysicalDeviceVariablePointersFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceVariablePointersFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    variable_pointers_storage_buffer Bool32
    variable_pointers      Bool32
} 

pub type PhysicalDeviceVariablePointerFeatures = PhysicalDeviceVariablePointersFeatures

// PhysicalDeviceProtectedMemoryFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceProtectedMemoryFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    protected_memory       Bool32
} 

// PhysicalDeviceProtectedMemoryProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceProtectedMemoryProperties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    protected_no_fault     Bool32
} 

pub struct DeviceQueueInfo2 {
mut:
    s_type                          StructureType
    p_next                          voidptr
    flags                           DeviceQueueCreateFlags
    queue_family_index              u32
    queue_index                     u32
} 

// ProtectedSubmitInfo extends VkSubmitInfo
pub struct ProtectedSubmitInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    protected_submit       Bool32
} 

pub struct SamplerYcbcrConversionCreateInfo {
mut:
    s_type                               StructureType
    p_next                               voidptr
    format                               Format
    ycbcr_model                          SamplerYcbcrModelConversion
    ycbcr_range                          SamplerYcbcrRange
    components                           ComponentMapping
    x_chroma_offset                      ChromaLocation
    y_chroma_offset                      ChromaLocation
    chroma_filter                        Filter
    force_explicit_reconstruction        Bool32
} 

// SamplerYcbcrConversionInfo extends VkSamplerCreateInfo,VkImageViewCreateInfo
pub struct SamplerYcbcrConversionInfo {
mut:
    s_type                          StructureType
    p_next                          voidptr
    conversion                      C.SamplerYcbcrConversion
} 

// BindImagePlaneMemoryInfo extends VkBindImageMemoryInfo
pub struct BindImagePlaneMemoryInfo {
mut:
    s_type                       StructureType
    p_next                       voidptr
    plane_aspect                 ImageAspectFlagBits
} 

// ImagePlaneMemoryRequirementsInfo extends VkImageMemoryRequirementsInfo2
pub struct ImagePlaneMemoryRequirementsInfo {
mut:
    s_type                       StructureType
    p_next                       voidptr
    plane_aspect                 ImageAspectFlagBits
} 

// PhysicalDeviceSamplerYcbcrConversionFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceSamplerYcbcrConversionFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    sampler_ycbcr_conversion Bool32
} 

// SamplerYcbcrConversionImageFormatProperties extends VkImageFormatProperties2
pub struct SamplerYcbcrConversionImageFormatProperties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    combined_image_sampler_descriptor_count u32
} 

pub struct DescriptorUpdateTemplateEntry {
mut:
    dst_binding             u32
    dst_array_element       u32
    descriptor_count        u32
    descriptor_type         DescriptorType
    offset                  usize
    stride                  usize
} 

pub struct DescriptorUpdateTemplateCreateInfo {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    flags                                         DescriptorUpdateTemplateCreateFlags
    descriptor_update_entry_count                 u32
    p_descriptor_update_entries                   &DescriptorUpdateTemplateEntry
    template_type                                 DescriptorUpdateTemplateType
    descriptor_set_layout                         C.DescriptorSetLayout
    pipeline_bind_point                           PipelineBindPoint
    pipeline_layout                               C.PipelineLayout
    set                                           u32
} 

pub struct ExternalMemoryProperties {
mut:
    external_memory_features               ExternalMemoryFeatureFlags
    export_from_imported_handle_types      ExternalMemoryHandleTypeFlags
    compatible_handle_types                ExternalMemoryHandleTypeFlags
} 

// PhysicalDeviceExternalImageFormatInfo extends VkPhysicalDeviceImageFormatInfo2
pub struct PhysicalDeviceExternalImageFormatInfo {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    handle_type                               ExternalMemoryHandleTypeFlagBits
} 

// ExternalImageFormatProperties extends VkImageFormatProperties2
pub struct ExternalImageFormatProperties {
mut:
    s_type                            StructureType
    p_next                            voidptr
    external_memory_properties        ExternalMemoryProperties
} 

pub struct PhysicalDeviceExternalBufferInfo {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    flags                                     BufferCreateFlags
    usage                                     BufferUsageFlags
    handle_type                               ExternalMemoryHandleTypeFlagBits
} 

pub struct ExternalBufferProperties {
mut:
    s_type                            StructureType
    p_next                            voidptr
    external_memory_properties        ExternalMemoryProperties
} 

// PhysicalDeviceIDProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceIDProperties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_uuid            []u8
    driver_uuid            []u8
    device_luid            []u8
    device_node_mask       u32
    device_luid_valid      Bool32
} 

// ExternalMemoryImageCreateInfo extends VkImageCreateInfo
pub struct ExternalMemoryImageCreateInfo {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    handle_types                           ExternalMemoryHandleTypeFlags
} 

// ExternalMemoryBufferCreateInfo extends VkBufferCreateInfo
pub struct ExternalMemoryBufferCreateInfo {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    handle_types                           ExternalMemoryHandleTypeFlags
} 

// ExportMemoryAllocateInfo extends VkMemoryAllocateInfo
pub struct ExportMemoryAllocateInfo {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    handle_types                           ExternalMemoryHandleTypeFlags
} 

pub struct PhysicalDeviceExternalFenceInfo {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    handle_type                              ExternalFenceHandleTypeFlagBits
} 

pub struct ExternalFenceProperties {
mut:
    s_type                                StructureType
    p_next                                voidptr
    export_from_imported_handle_types     ExternalFenceHandleTypeFlags
    compatible_handle_types               ExternalFenceHandleTypeFlags
    external_fence_features               ExternalFenceFeatureFlags
} 

// ExportFenceCreateInfo extends VkFenceCreateInfo
pub struct ExportFenceCreateInfo {
mut:
    s_type                                StructureType
    p_next                                voidptr
    handle_types                          ExternalFenceHandleTypeFlags
} 

// ExportSemaphoreCreateInfo extends VkSemaphoreCreateInfo
pub struct ExportSemaphoreCreateInfo {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    handle_types                              ExternalSemaphoreHandleTypeFlags
} 

pub struct PhysicalDeviceExternalSemaphoreInfo {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    handle_type                                  ExternalSemaphoreHandleTypeFlagBits
} 

pub struct ExternalSemaphoreProperties {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    export_from_imported_handle_types         ExternalSemaphoreHandleTypeFlags
    compatible_handle_types                   ExternalSemaphoreHandleTypeFlags
    external_semaphore_features               ExternalSemaphoreFeatureFlags
} 

// PhysicalDeviceMaintenance3Properties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceMaintenance3Properties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_per_set_descriptors u32
    max_memory_allocation_size DeviceSize
} 

pub struct DescriptorSetLayoutSupport {
mut:
    s_type                 StructureType
    p_next                 voidptr
    supported              Bool32
} 

// PhysicalDeviceShaderDrawParametersFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderDrawParametersFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_draw_parameters Bool32
} 

pub type PhysicalDeviceShaderDrawParameterFeatures = PhysicalDeviceShaderDrawParametersFeatures

type VkEnumerateInstanceVersion = fn (     &u32) Result

pub fn enumerate_instance_version(
    p_api_version                                   &u32) Result {
      f := VkEnumerateInstanceVersion((*loader_p).get_sym('vkEnumerateInstanceVersion'
    ) or { 
        println("Couldn't load symbol for 'vkEnumerateInstanceVersion': ${err}")
        return Result.error_unknown
    })
    return f(
    p_api_version)
}


type VkBindBufferMemory2 = fn (     C.Device,     u32,     &BindBufferMemoryInfo) Result

pub fn bind_buffer_memory2(
    device                                          C.Device,
    bind_info_count                                 u32,
    p_bind_infos                                    &BindBufferMemoryInfo) Result {
      f := VkBindBufferMemory2((*loader_p).get_sym('vkBindBufferMemory2'
    ) or { 
        println("Couldn't load symbol for 'vkBindBufferMemory2': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    bind_info_count,
    p_bind_infos)
}


type VkBindImageMemory2 = fn (     C.Device,     u32,     &BindImageMemoryInfo) Result

pub fn bind_image_memory2(
    device                                          C.Device,
    bind_info_count                                 u32,
    p_bind_infos                                    &BindImageMemoryInfo) Result {
      f := VkBindImageMemory2((*loader_p).get_sym('vkBindImageMemory2'
    ) or { 
        println("Couldn't load symbol for 'vkBindImageMemory2': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    bind_info_count,
    p_bind_infos)
}


type VkGetDeviceGroupPeerMemoryFeatures = fn (     C.Device,     u32,     u32,     u32,     &PeerMemoryFeatureFlags) 

pub fn get_device_group_peer_memory_features(
    device                                          C.Device,
    heap_index                                      u32,
    local_device_index                              u32,
    remote_device_index                             u32,
    p_peer_memory_features                          &PeerMemoryFeatureFlags)  {
      f := VkGetDeviceGroupPeerMemoryFeatures((*loader_p).get_sym('vkGetDeviceGroupPeerMemoryFeatures'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceGroupPeerMemoryFeatures': ${err}")
        return 
    })
    f(
    device,
    heap_index,
    local_device_index,
    remote_device_index,
    p_peer_memory_features)
}


type VkCmdSetDeviceMask = fn (     C.CommandBuffer,     u32) 

pub fn cmd_set_device_mask(
    command_buffer                                  C.CommandBuffer,
    device_mask                                     u32)  {
      f := VkCmdSetDeviceMask((*loader_p).get_sym('vkCmdSetDeviceMask'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDeviceMask': ${err}")
        return 
    })
    f(
    command_buffer,
    device_mask)
}


type VkCmdDispatchBase = fn (     C.CommandBuffer,     u32,     u32,     u32,     u32,     u32,     u32) 

pub fn cmd_dispatch_base(
    command_buffer                                  C.CommandBuffer,
    base_group_x                                    u32,
    base_group_y                                    u32,
    base_group_z                                    u32,
    group_count_x                                   u32,
    group_count_y                                   u32,
    group_count_z                                   u32)  {
      f := VkCmdDispatchBase((*loader_p).get_sym('vkCmdDispatchBase'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDispatchBase': ${err}")
        return 
    })
    f(
    command_buffer,
    base_group_x,
    base_group_y,
    base_group_z,
    group_count_x,
    group_count_y,
    group_count_z)
}


type VkEnumeratePhysicalDeviceGroups = fn (     C.Instance,     &u32,     &PhysicalDeviceGroupProperties) Result

pub fn enumerate_physical_device_groups(
    instance                                        C.Instance,
    p_physical_device_group_count                   &u32,
    p_physical_device_group_properties              &PhysicalDeviceGroupProperties) Result {
      f := VkEnumeratePhysicalDeviceGroups((*loader_p).get_sym('vkEnumeratePhysicalDeviceGroups'
    ) or { 
        println("Couldn't load symbol for 'vkEnumeratePhysicalDeviceGroups': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_physical_device_group_count,
    p_physical_device_group_properties)
}


type VkGetImageMemoryRequirements2 = fn (     C.Device,     &ImageMemoryRequirementsInfo2,     &MemoryRequirements2) 

pub fn get_image_memory_requirements2(
    device                                          C.Device,
    p_info                                          &ImageMemoryRequirementsInfo2,
    p_memory_requirements                           &MemoryRequirements2)  {
      f := VkGetImageMemoryRequirements2((*loader_p).get_sym('vkGetImageMemoryRequirements2'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageMemoryRequirements2': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_memory_requirements)
}


type VkGetBufferMemoryRequirements2 = fn (     C.Device,     &BufferMemoryRequirementsInfo2,     &MemoryRequirements2) 

pub fn get_buffer_memory_requirements2(
    device                                          C.Device,
    p_info                                          &BufferMemoryRequirementsInfo2,
    p_memory_requirements                           &MemoryRequirements2)  {
      f := VkGetBufferMemoryRequirements2((*loader_p).get_sym('vkGetBufferMemoryRequirements2'
    ) or { 
        println("Couldn't load symbol for 'vkGetBufferMemoryRequirements2': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_memory_requirements)
}


type VkGetImageSparseMemoryRequirements2 = fn (     C.Device,     &ImageSparseMemoryRequirementsInfo2,     &u32,     &SparseImageMemoryRequirements2) 

pub fn get_image_sparse_memory_requirements2(
    device                                          C.Device,
    p_info                                          &ImageSparseMemoryRequirementsInfo2,
    p_sparse_memory_requirement_count               &u32,
    p_sparse_memory_requirements                    &SparseImageMemoryRequirements2)  {
      f := VkGetImageSparseMemoryRequirements2((*loader_p).get_sym('vkGetImageSparseMemoryRequirements2'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageSparseMemoryRequirements2': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_sparse_memory_requirement_count,
    p_sparse_memory_requirements)
}


type VkGetPhysicalDeviceFeatures2 = fn (     C.PhysicalDevice,     &PhysicalDeviceFeatures2) 

pub fn get_physical_device_features2(
    physical_device                                 C.PhysicalDevice,
    p_features                                      &PhysicalDeviceFeatures2)  {
      f := VkGetPhysicalDeviceFeatures2((*loader_p).get_sym('vkGetPhysicalDeviceFeatures2'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceFeatures2': ${err}")
        return 
    })
    f(
    physical_device,
    p_features)
}


type VkGetPhysicalDeviceProperties2 = fn (     C.PhysicalDevice,     &PhysicalDeviceProperties2) 

pub fn get_physical_device_properties2(
    physical_device                                 C.PhysicalDevice,
    p_properties                                    &PhysicalDeviceProperties2)  {
      f := VkGetPhysicalDeviceProperties2((*loader_p).get_sym('vkGetPhysicalDeviceProperties2'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceProperties2': ${err}")
        return 
    })
    f(
    physical_device,
    p_properties)
}


type VkGetPhysicalDeviceFormatProperties2 = fn (     C.PhysicalDevice,     Format,     &FormatProperties2) 

pub fn get_physical_device_format_properties2(
    physical_device                                 C.PhysicalDevice,
    format                                          Format,
    p_format_properties                             &FormatProperties2)  {
      f := VkGetPhysicalDeviceFormatProperties2((*loader_p).get_sym('vkGetPhysicalDeviceFormatProperties2'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceFormatProperties2': ${err}")
        return 
    })
    f(
    physical_device,
    format,
    p_format_properties)
}


type VkGetPhysicalDeviceImageFormatProperties2 = fn (     C.PhysicalDevice,     &PhysicalDeviceImageFormatInfo2,     &ImageFormatProperties2) Result

pub fn get_physical_device_image_format_properties2(
    physical_device                                 C.PhysicalDevice,
    p_image_format_info                             &PhysicalDeviceImageFormatInfo2,
    p_image_format_properties                       &ImageFormatProperties2) Result {
      f := VkGetPhysicalDeviceImageFormatProperties2((*loader_p).get_sym('vkGetPhysicalDeviceImageFormatProperties2'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceImageFormatProperties2': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_image_format_info,
    p_image_format_properties)
}


type VkGetPhysicalDeviceQueueFamilyProperties2 = fn (     C.PhysicalDevice,     &u32,     &QueueFamilyProperties2) 

pub fn get_physical_device_queue_family_properties2(
    physical_device                                 C.PhysicalDevice,
    p_queue_family_property_count                   &u32,
    p_queue_family_properties                       &QueueFamilyProperties2)  {
      f := VkGetPhysicalDeviceQueueFamilyProperties2((*loader_p).get_sym('vkGetPhysicalDeviceQueueFamilyProperties2'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceQueueFamilyProperties2': ${err}")
        return 
    })
    f(
    physical_device,
    p_queue_family_property_count,
    p_queue_family_properties)
}


type VkGetPhysicalDeviceMemoryProperties2 = fn (     C.PhysicalDevice,     &PhysicalDeviceMemoryProperties2) 

pub fn get_physical_device_memory_properties2(
    physical_device                                 C.PhysicalDevice,
    p_memory_properties                             &PhysicalDeviceMemoryProperties2)  {
      f := VkGetPhysicalDeviceMemoryProperties2((*loader_p).get_sym('vkGetPhysicalDeviceMemoryProperties2'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceMemoryProperties2': ${err}")
        return 
    })
    f(
    physical_device,
    p_memory_properties)
}


type VkGetPhysicalDeviceSparseImageFormatProperties2 = fn (     C.PhysicalDevice,     &PhysicalDeviceSparseImageFormatInfo2,     &u32,     &SparseImageFormatProperties2) 

pub fn get_physical_device_sparse_image_format_properties2(
    physical_device                                 C.PhysicalDevice,
    p_format_info                                   &PhysicalDeviceSparseImageFormatInfo2,
    p_property_count                                &u32,
    p_properties                                    &SparseImageFormatProperties2)  {
      f := VkGetPhysicalDeviceSparseImageFormatProperties2((*loader_p).get_sym('vkGetPhysicalDeviceSparseImageFormatProperties2'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSparseImageFormatProperties2': ${err}")
        return 
    })
    f(
    physical_device,
    p_format_info,
    p_property_count,
    p_properties)
}


type VkTrimCommandPool = fn (     C.Device,     C.CommandPool,     CommandPoolTrimFlags) 

pub fn trim_command_pool(
    device                                          C.Device,
    command_pool                                    C.CommandPool,
    flags                                           CommandPoolTrimFlags)  {
      f := VkTrimCommandPool((*loader_p).get_sym('vkTrimCommandPool'
    ) or { 
        println("Couldn't load symbol for 'vkTrimCommandPool': ${err}")
        return 
    })
    f(
    device,
    command_pool,
    flags)
}


type VkGetDeviceQueue2 = fn (     C.Device,     &DeviceQueueInfo2,     &C.Queue) 

pub fn get_device_queue2(
    device                                          C.Device,
    p_queue_info                                    &DeviceQueueInfo2,
    p_queue                                         &C.Queue)  {
      f := VkGetDeviceQueue2((*loader_p).get_sym('vkGetDeviceQueue2'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceQueue2': ${err}")
        return 
    })
    f(
    device,
    p_queue_info,
    p_queue)
}


type VkCreateSamplerYcbcrConversion = fn (     C.Device,     &SamplerYcbcrConversionCreateInfo,     &AllocationCallbacks,     &C.SamplerYcbcrConversion) Result

pub fn create_sampler_ycbcr_conversion(
    device                                          C.Device,
    p_create_info                                   &SamplerYcbcrConversionCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_ycbcr_conversion                              &C.SamplerYcbcrConversion) Result {
      f := VkCreateSamplerYcbcrConversion((*loader_p).get_sym('vkCreateSamplerYcbcrConversion'
    ) or { 
        println("Couldn't load symbol for 'vkCreateSamplerYcbcrConversion': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_ycbcr_conversion)
}


type VkDestroySamplerYcbcrConversion = fn (     C.Device,     C.SamplerYcbcrConversion,     &AllocationCallbacks) 

pub fn destroy_sampler_ycbcr_conversion(
    device                                          C.Device,
    ycbcr_conversion                                C.SamplerYcbcrConversion,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroySamplerYcbcrConversion((*loader_p).get_sym('vkDestroySamplerYcbcrConversion'
    ) or { 
        println("Couldn't load symbol for 'vkDestroySamplerYcbcrConversion': ${err}")
        return 
    })
    f(
    device,
    ycbcr_conversion,
    p_allocator)
}


type VkCreateDescriptorUpdateTemplate = fn (     C.Device,     &DescriptorUpdateTemplateCreateInfo,     &AllocationCallbacks,     &C.DescriptorUpdateTemplate) Result

pub fn create_descriptor_update_template(
    device                                          C.Device,
    p_create_info                                   &DescriptorUpdateTemplateCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_descriptor_update_template                    &C.DescriptorUpdateTemplate) Result {
      f := VkCreateDescriptorUpdateTemplate((*loader_p).get_sym('vkCreateDescriptorUpdateTemplate'
    ) or { 
        println("Couldn't load symbol for 'vkCreateDescriptorUpdateTemplate': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_descriptor_update_template)
}


type VkDestroyDescriptorUpdateTemplate = fn (     C.Device,     C.DescriptorUpdateTemplate,     &AllocationCallbacks) 

pub fn destroy_descriptor_update_template(
    device                                          C.Device,
    descriptor_update_template                      C.DescriptorUpdateTemplate,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyDescriptorUpdateTemplate((*loader_p).get_sym('vkDestroyDescriptorUpdateTemplate'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyDescriptorUpdateTemplate': ${err}")
        return 
    })
    f(
    device,
    descriptor_update_template,
    p_allocator)
}


type VkUpdateDescriptorSetWithTemplate = fn (     C.Device,     C.DescriptorSet,     C.DescriptorUpdateTemplate,     voidptr) 

pub fn update_descriptor_set_with_template(
    device                                          C.Device,
    descriptor_set                                  C.DescriptorSet,
    descriptor_update_template                      C.DescriptorUpdateTemplate,
    p_data                                          voidptr)  {
      f := VkUpdateDescriptorSetWithTemplate((*loader_p).get_sym('vkUpdateDescriptorSetWithTemplate'
    ) or { 
        println("Couldn't load symbol for 'vkUpdateDescriptorSetWithTemplate': ${err}")
        return 
    })
    f(
    device,
    descriptor_set,
    descriptor_update_template,
    p_data)
}


type VkGetPhysicalDeviceExternalBufferProperties = fn (     C.PhysicalDevice,     &PhysicalDeviceExternalBufferInfo,     &ExternalBufferProperties) 

pub fn get_physical_device_external_buffer_properties(
    physical_device                                 C.PhysicalDevice,
    p_external_buffer_info                          &PhysicalDeviceExternalBufferInfo,
    p_external_buffer_properties                    &ExternalBufferProperties)  {
      f := VkGetPhysicalDeviceExternalBufferProperties((*loader_p).get_sym('vkGetPhysicalDeviceExternalBufferProperties'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceExternalBufferProperties': ${err}")
        return 
    })
    f(
    physical_device,
    p_external_buffer_info,
    p_external_buffer_properties)
}


type VkGetPhysicalDeviceExternalFenceProperties = fn (     C.PhysicalDevice,     &PhysicalDeviceExternalFenceInfo,     &ExternalFenceProperties) 

pub fn get_physical_device_external_fence_properties(
    physical_device                                 C.PhysicalDevice,
    p_external_fence_info                           &PhysicalDeviceExternalFenceInfo,
    p_external_fence_properties                     &ExternalFenceProperties)  {
      f := VkGetPhysicalDeviceExternalFenceProperties((*loader_p).get_sym('vkGetPhysicalDeviceExternalFenceProperties'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceExternalFenceProperties': ${err}")
        return 
    })
    f(
    physical_device,
    p_external_fence_info,
    p_external_fence_properties)
}


type VkGetPhysicalDeviceExternalSemaphoreProperties = fn (     C.PhysicalDevice,     &PhysicalDeviceExternalSemaphoreInfo,     &ExternalSemaphoreProperties) 

pub fn get_physical_device_external_semaphore_properties(
    physical_device                                 C.PhysicalDevice,
    p_external_semaphore_info                       &PhysicalDeviceExternalSemaphoreInfo,
    p_external_semaphore_properties                 &ExternalSemaphoreProperties)  {
      f := VkGetPhysicalDeviceExternalSemaphoreProperties((*loader_p).get_sym('vkGetPhysicalDeviceExternalSemaphoreProperties'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceExternalSemaphoreProperties': ${err}")
        return 
    })
    f(
    physical_device,
    p_external_semaphore_info,
    p_external_semaphore_properties)
}


type VkGetDescriptorSetLayoutSupport = fn (     C.Device,     &DescriptorSetLayoutCreateInfo,     &DescriptorSetLayoutSupport) 

pub fn get_descriptor_set_layout_support(
    device                                          C.Device,
    p_create_info                                   &DescriptorSetLayoutCreateInfo,
    p_support                                       &DescriptorSetLayoutSupport)  {
      f := VkGetDescriptorSetLayoutSupport((*loader_p).get_sym('vkGetDescriptorSetLayoutSupport'
    ) or { 
        println("Couldn't load symbol for 'vkGetDescriptorSetLayoutSupport': ${err}")
        return 
    })
    f(
    device,
    p_create_info,
    p_support)
}




// VK_VERSION_1_2 is a preprocessor guard. Do not pass it to API calls.
const version_1_2 = 1
// Vulkan 1.2 version number
pub const api_version_1_2 = make_api_version(0, 1, 2, 0)// Patch version should always be set to 0

pub const max_driver_name_size              = u32(256)
pub const max_driver_info_size              = u32(256)

pub enum DriverId {
    driver_id_amd_proprietary = int(1)
    driver_id_amd_open_source = int(2)
    driver_id_mesa_radv = int(3)
    driver_id_nvidia_proprietary = int(4)
    driver_id_intel_proprietary_windows = int(5)
    driver_id_intel_open_source_mesa = int(6)
    driver_id_imagination_proprietary = int(7)
    driver_id_qualcomm_proprietary = int(8)
    driver_id_arm_proprietary = int(9)
    driver_id_google_swiftshader = int(10)
    driver_id_ggp_proprietary = int(11)
    driver_id_broadcom_proprietary = int(12)
    driver_id_mesa_llvmpipe = int(13)
    driver_id_moltenvk = int(14)
    driver_id_coreavi_proprietary = int(15)
    driver_id_juice_proprietary = int(16)
    driver_id_verisilicon_proprietary = int(17)
    driver_id_mesa_turnip = int(18)
    driver_id_mesa_v3dv = int(19)
    driver_id_mesa_panvk = int(20)
    driver_id_samsung_proprietary = int(21)
    driver_id_mesa_venus = int(22)
    driver_id_mesa_dozen = int(23)
    driver_id_mesa_nvk = int(24)
    driver_id_imagination_open_source_mesa = int(25)
    driver_id_mesa_agxv = int(26)
    driver_id_max_enum = int(0x7FFFFFFF)
}


pub enum ShaderFloatControlsIndependence {
    shader_float_controls_independence_32_bit_only = int(0)
    shader_float_controls_independence_all = int(1)
    shader_float_controls_independence_none = int(2)
    shader_float_controls_independence_max_enum = int(0x7FFFFFFF)
}


pub enum SamplerReductionMode {
    sampler_reduction_mode_weighted_average = int(0)
    sampler_reduction_mode_min = int(1)
    sampler_reduction_mode_max = int(2)
    sampler_reduction_mode_weighted_average_rangeclamp_qcom = int(1000521000)
    sampler_reduction_mode_max_enum = int(0x7FFFFFFF)
}


pub enum SemaphoreType {
    semaphore_type_binary = int(0)
    semaphore_type_timeline = int(1)
    semaphore_type_max_enum = int(0x7FFFFFFF)
}


pub enum ResolveModeFlagBits {
    resolve_mode_none = int(0)
    resolve_mode_sample_zero_bit = int(0x00000001)
    resolve_mode_average_bit = int(0x00000002)
    resolve_mode_min_bit = int(0x00000004)
    resolve_mode_max_bit = int(0x00000008)
    resolve_mode_external_format_downsample_android = int(0x00000010)
    resolve_mode_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ResolveModeFlags = u32

pub enum DescriptorBindingFlagBits {
    descriptor_binding_update_after_bind_bit = int(0x00000001)
    descriptor_binding_update_unused_while_pending_bit = int(0x00000002)
    descriptor_binding_partially_bound_bit = int(0x00000004)
    descriptor_binding_variable_descriptor_count_bit = int(0x00000008)
    descriptor_binding_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type DescriptorBindingFlags = u32

pub enum SemaphoreWaitFlagBits {
    semaphore_wait_any_bit = int(0x00000001)
    semaphore_wait_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type SemaphoreWaitFlags = u32
// PhysicalDeviceVulkan11Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceVulkan11Features {
mut:
    s_type                 StructureType
    p_next                 voidptr
    storage_buffer16_bit_access Bool32
    uniform_and_storage_buffer16_bit_access Bool32
    storage_push_constant16 Bool32
    storage_input_output16 Bool32
    multiview              Bool32
    multiview_geometry_shader Bool32
    multiview_tessellation_shader Bool32
    variable_pointers_storage_buffer Bool32
    variable_pointers      Bool32
    protected_memory       Bool32
    sampler_ycbcr_conversion Bool32
    shader_draw_parameters Bool32
} 

// PhysicalDeviceVulkan11Properties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceVulkan11Properties {
mut:
    s_type                         StructureType
    p_next                         voidptr
    device_uuid                    []u8
    driver_uuid                    []u8
    device_luid                    []u8
    device_node_mask               u32
    device_luid_valid              Bool32
    subgroup_size                  u32
    subgroup_supported_stages      ShaderStageFlags
    subgroup_supported_operations  SubgroupFeatureFlags
    subgroup_quad_operations_in_all_stages Bool32
    point_clipping_behavior        PointClippingBehavior
    max_multiview_view_count       u32
    max_multiview_instance_index   u32
    protected_no_fault             Bool32
    max_per_set_descriptors        u32
    max_memory_allocation_size     DeviceSize
} 

// PhysicalDeviceVulkan12Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceVulkan12Features {
mut:
    s_type                 StructureType
    p_next                 voidptr
    sampler_mirror_clamp_to_edge Bool32
    draw_indirect_count    Bool32
    storage_buffer8_bit_access Bool32
    uniform_and_storage_buffer8_bit_access Bool32
    storage_push_constant8 Bool32
    shader_buffer_int64_atomics Bool32
    shader_shared_int64_atomics Bool32
    shader_float16         Bool32
    shader_int8            Bool32
    descriptor_indexing    Bool32
    shader_input_attachment_array_dynamic_indexing Bool32
    shader_uniform_texel_buffer_array_dynamic_indexing Bool32
    shader_storage_texel_buffer_array_dynamic_indexing Bool32
    shader_uniform_buffer_array_non_uniform_indexing Bool32
    shader_sampled_image_array_non_uniform_indexing Bool32
    shader_storage_buffer_array_non_uniform_indexing Bool32
    shader_storage_image_array_non_uniform_indexing Bool32
    shader_input_attachment_array_non_uniform_indexing Bool32
    shader_uniform_texel_buffer_array_non_uniform_indexing Bool32
    shader_storage_texel_buffer_array_non_uniform_indexing Bool32
    descriptor_binding_uniform_buffer_update_after_bind Bool32
    descriptor_binding_sampled_image_update_after_bind Bool32
    descriptor_binding_storage_image_update_after_bind Bool32
    descriptor_binding_storage_buffer_update_after_bind Bool32
    descriptor_binding_uniform_texel_buffer_update_after_bind Bool32
    descriptor_binding_storage_texel_buffer_update_after_bind Bool32
    descriptor_binding_update_unused_while_pending Bool32
    descriptor_binding_partially_bound Bool32
    descriptor_binding_variable_descriptor_count Bool32
    runtime_descriptor_array Bool32
    sampler_filter_minmax  Bool32
    scalar_block_layout    Bool32
    imageless_framebuffer  Bool32
    uniform_buffer_standard_layout Bool32
    shader_subgroup_extended_types Bool32
    separate_depth_stencil_layouts Bool32
    host_query_reset       Bool32
    timeline_semaphore     Bool32
    buffer_device_address  Bool32
    buffer_device_address_capture_replay Bool32
    buffer_device_address_multi_device Bool32
    vulkan_memory_model    Bool32
    vulkan_memory_model_device_scope Bool32
    vulkan_memory_model_availability_visibility_chains Bool32
    shader_output_viewport_index Bool32
    shader_output_layer    Bool32
    subgroup_broadcast_dynamic_id Bool32
} 

pub struct ConformanceVersion {
mut:
    major          u8
    minor          u8
    subminor       u8
    patch          u8
} 

// PhysicalDeviceVulkan12Properties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceVulkan12Properties {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    driver_id                                DriverId
    driver_name                              []char
    driver_info                              []char
    conformance_version                      ConformanceVersion
    denorm_behavior_independence             ShaderFloatControlsIndependence
    rounding_mode_independence               ShaderFloatControlsIndependence
    shader_signed_zero_inf_nan_preserve_float16 Bool32
    shader_signed_zero_inf_nan_preserve_float32 Bool32
    shader_signed_zero_inf_nan_preserve_float64 Bool32
    shader_denorm_preserve_float16           Bool32
    shader_denorm_preserve_float32           Bool32
    shader_denorm_preserve_float64           Bool32
    shader_denorm_flush_to_zero_float16      Bool32
    shader_denorm_flush_to_zero_float32      Bool32
    shader_denorm_flush_to_zero_float64      Bool32
    shader_rounding_mode_rte_float16         Bool32
    shader_rounding_mode_rte_float32         Bool32
    shader_rounding_mode_rte_float64         Bool32
    shader_rounding_mode_rtz_float16         Bool32
    shader_rounding_mode_rtz_float32         Bool32
    shader_rounding_mode_rtz_float64         Bool32
    max_update_after_bind_descriptors_in_all_pools u32
    shader_uniform_buffer_array_non_uniform_indexing_native Bool32
    shader_sampled_image_array_non_uniform_indexing_native Bool32
    shader_storage_buffer_array_non_uniform_indexing_native Bool32
    shader_storage_image_array_non_uniform_indexing_native Bool32
    shader_input_attachment_array_non_uniform_indexing_native Bool32
    robust_buffer_access_update_after_bind   Bool32
    quad_divergent_implicit_lod              Bool32
    max_per_stage_descriptor_update_after_bind_samplers u32
    max_per_stage_descriptor_update_after_bind_uniform_buffers u32
    max_per_stage_descriptor_update_after_bind_storage_buffers u32
    max_per_stage_descriptor_update_after_bind_sampled_images u32
    max_per_stage_descriptor_update_after_bind_storage_images u32
    max_per_stage_descriptor_update_after_bind_input_attachments u32
    max_per_stage_update_after_bind_resources u32
    max_descriptor_set_update_after_bind_samplers u32
    max_descriptor_set_update_after_bind_uniform_buffers u32
    max_descriptor_set_update_after_bind_uniform_buffers_dynamic u32
    max_descriptor_set_update_after_bind_storage_buffers u32
    max_descriptor_set_update_after_bind_storage_buffers_dynamic u32
    max_descriptor_set_update_after_bind_sampled_images u32
    max_descriptor_set_update_after_bind_storage_images u32
    max_descriptor_set_update_after_bind_input_attachments u32
    supported_depth_resolve_modes            ResolveModeFlags
    supported_stencil_resolve_modes          ResolveModeFlags
    independent_resolve_none                 Bool32
    independent_resolve                      Bool32
    filter_minmax_single_component_formats   Bool32
    filter_minmax_image_component_mapping    Bool32
    max_timeline_semaphore_value_difference  u64
    framebuffer_integer_color_sample_counts  SampleCountFlags
} 

// ImageFormatListCreateInfo extends VkImageCreateInfo,VkSwapchainCreateInfoKHR,VkPhysicalDeviceImageFormatInfo2
pub struct ImageFormatListCreateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    view_format_count      u32
    p_view_formats         &Format
} 

pub struct AttachmentDescription2 {
mut:
    s_type                              StructureType
    p_next                              voidptr
    flags                               AttachmentDescriptionFlags
    format                              Format
    samples                             SampleCountFlagBits
    load_op                             AttachmentLoadOp
    store_op                            AttachmentStoreOp
    stencil_load_op                     AttachmentLoadOp
    stencil_store_op                    AttachmentStoreOp
    initial_layout                      ImageLayout
    final_layout                        ImageLayout
} 

pub struct AttachmentReference2 {
mut:
    s_type                    StructureType
    p_next                    voidptr
    attachment                u32
    layout                    ImageLayout
    aspect_mask               ImageAspectFlags
} 

pub struct SubpassDescription2 {
mut:
    s_type                               StructureType
    p_next                               voidptr
    flags                                SubpassDescriptionFlags
    pipeline_bind_point                  PipelineBindPoint
    view_mask                            u32
    input_attachment_count               u32
    p_input_attachments                  &AttachmentReference2
    color_attachment_count               u32
    p_color_attachments                  &AttachmentReference2
    p_resolve_attachments                &AttachmentReference2
    p_depth_stencil_attachment           &AttachmentReference2
    preserve_attachment_count            u32
    p_preserve_attachments               &u32
} 

pub struct SubpassDependency2 {
mut:
    s_type                      StructureType
    p_next                      voidptr
    src_subpass                 u32
    dst_subpass                 u32
    src_stage_mask              PipelineStageFlags
    dst_stage_mask              PipelineStageFlags
    src_access_mask             AccessFlags
    dst_access_mask             AccessFlags
    dependency_flags            DependencyFlags
    view_offset                 i32
} 

pub struct RenderPassCreateInfo2 {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    flags                                  RenderPassCreateFlags
    attachment_count                       u32
    p_attachments                          &AttachmentDescription2
    subpass_count                          u32
    p_subpasses                            &SubpassDescription2
    dependency_count                       u32
    p_dependencies                         &SubpassDependency2
    correlated_view_mask_count             u32
    p_correlated_view_masks                &u32
} 

pub struct SubpassBeginInfo {
mut:
    s_type                   StructureType
    p_next                   voidptr
    contents                 SubpassContents
} 

pub struct SubpassEndInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
} 

// PhysicalDevice8BitStorageFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevice8BitStorageFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    storage_buffer8_bit_access Bool32
    uniform_and_storage_buffer8_bit_access Bool32
    storage_push_constant8 Bool32
} 

// PhysicalDeviceDriverProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceDriverProperties {
mut:
    s_type                      StructureType
    p_next                      voidptr
    driver_id                   DriverId
    driver_name                 []char
    driver_info                 []char
    conformance_version         ConformanceVersion
} 

// PhysicalDeviceShaderAtomicInt64Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderAtomicInt64Features {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_buffer_int64_atomics Bool32
    shader_shared_int64_atomics Bool32
} 

// PhysicalDeviceShaderFloat16Int8Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderFloat16Int8Features {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_float16         Bool32
    shader_int8            Bool32
} 

// PhysicalDeviceFloatControlsProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceFloatControlsProperties {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    denorm_behavior_independence             ShaderFloatControlsIndependence
    rounding_mode_independence               ShaderFloatControlsIndependence
    shader_signed_zero_inf_nan_preserve_float16 Bool32
    shader_signed_zero_inf_nan_preserve_float32 Bool32
    shader_signed_zero_inf_nan_preserve_float64 Bool32
    shader_denorm_preserve_float16           Bool32
    shader_denorm_preserve_float32           Bool32
    shader_denorm_preserve_float64           Bool32
    shader_denorm_flush_to_zero_float16      Bool32
    shader_denorm_flush_to_zero_float32      Bool32
    shader_denorm_flush_to_zero_float64      Bool32
    shader_rounding_mode_rte_float16         Bool32
    shader_rounding_mode_rte_float32         Bool32
    shader_rounding_mode_rte_float64         Bool32
    shader_rounding_mode_rtz_float16         Bool32
    shader_rounding_mode_rtz_float32         Bool32
    shader_rounding_mode_rtz_float64         Bool32
} 

// DescriptorSetLayoutBindingFlagsCreateInfo extends VkDescriptorSetLayoutCreateInfo
pub struct DescriptorSetLayoutBindingFlagsCreateInfo {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    binding_count                          u32
    p_binding_flags                        &DescriptorBindingFlags
} 

// PhysicalDeviceDescriptorIndexingFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDescriptorIndexingFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_input_attachment_array_dynamic_indexing Bool32
    shader_uniform_texel_buffer_array_dynamic_indexing Bool32
    shader_storage_texel_buffer_array_dynamic_indexing Bool32
    shader_uniform_buffer_array_non_uniform_indexing Bool32
    shader_sampled_image_array_non_uniform_indexing Bool32
    shader_storage_buffer_array_non_uniform_indexing Bool32
    shader_storage_image_array_non_uniform_indexing Bool32
    shader_input_attachment_array_non_uniform_indexing Bool32
    shader_uniform_texel_buffer_array_non_uniform_indexing Bool32
    shader_storage_texel_buffer_array_non_uniform_indexing Bool32
    descriptor_binding_uniform_buffer_update_after_bind Bool32
    descriptor_binding_sampled_image_update_after_bind Bool32
    descriptor_binding_storage_image_update_after_bind Bool32
    descriptor_binding_storage_buffer_update_after_bind Bool32
    descriptor_binding_uniform_texel_buffer_update_after_bind Bool32
    descriptor_binding_storage_texel_buffer_update_after_bind Bool32
    descriptor_binding_update_unused_while_pending Bool32
    descriptor_binding_partially_bound Bool32
    descriptor_binding_variable_descriptor_count Bool32
    runtime_descriptor_array Bool32
} 

// PhysicalDeviceDescriptorIndexingProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceDescriptorIndexingProperties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_update_after_bind_descriptors_in_all_pools u32
    shader_uniform_buffer_array_non_uniform_indexing_native Bool32
    shader_sampled_image_array_non_uniform_indexing_native Bool32
    shader_storage_buffer_array_non_uniform_indexing_native Bool32
    shader_storage_image_array_non_uniform_indexing_native Bool32
    shader_input_attachment_array_non_uniform_indexing_native Bool32
    robust_buffer_access_update_after_bind Bool32
    quad_divergent_implicit_lod Bool32
    max_per_stage_descriptor_update_after_bind_samplers u32
    max_per_stage_descriptor_update_after_bind_uniform_buffers u32
    max_per_stage_descriptor_update_after_bind_storage_buffers u32
    max_per_stage_descriptor_update_after_bind_sampled_images u32
    max_per_stage_descriptor_update_after_bind_storage_images u32
    max_per_stage_descriptor_update_after_bind_input_attachments u32
    max_per_stage_update_after_bind_resources u32
    max_descriptor_set_update_after_bind_samplers u32
    max_descriptor_set_update_after_bind_uniform_buffers u32
    max_descriptor_set_update_after_bind_uniform_buffers_dynamic u32
    max_descriptor_set_update_after_bind_storage_buffers u32
    max_descriptor_set_update_after_bind_storage_buffers_dynamic u32
    max_descriptor_set_update_after_bind_sampled_images u32
    max_descriptor_set_update_after_bind_storage_images u32
    max_descriptor_set_update_after_bind_input_attachments u32
} 

// DescriptorSetVariableDescriptorCountAllocateInfo extends VkDescriptorSetAllocateInfo
pub struct DescriptorSetVariableDescriptorCountAllocateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    descriptor_set_count   u32
    p_descriptor_counts    &u32
} 

// DescriptorSetVariableDescriptorCountLayoutSupport extends VkDescriptorSetLayoutSupport
pub struct DescriptorSetVariableDescriptorCountLayoutSupport {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_variable_descriptor_count u32
} 

// SubpassDescriptionDepthStencilResolve extends VkSubpassDescription2
pub struct SubpassDescriptionDepthStencilResolve {
mut:
    s_type                               StructureType
    p_next                               voidptr
    depth_resolve_mode                   ResolveModeFlagBits
    stencil_resolve_mode                 ResolveModeFlagBits
    p_depth_stencil_resolve_attachment   &AttachmentReference2
} 

// PhysicalDeviceDepthStencilResolveProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceDepthStencilResolveProperties {
mut:
    s_type                    StructureType
    p_next                    voidptr
    supported_depth_resolve_modes ResolveModeFlags
    supported_stencil_resolve_modes ResolveModeFlags
    independent_resolve_none  Bool32
    independent_resolve       Bool32
} 

// PhysicalDeviceScalarBlockLayoutFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceScalarBlockLayoutFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    scalar_block_layout    Bool32
} 

// ImageStencilUsageCreateInfo extends VkImageCreateInfo,VkPhysicalDeviceImageFormatInfo2
pub struct ImageStencilUsageCreateInfo {
mut:
    s_type                   StructureType
    p_next                   voidptr
    stencil_usage            ImageUsageFlags
} 

// SamplerReductionModeCreateInfo extends VkSamplerCreateInfo
pub struct SamplerReductionModeCreateInfo {
mut:
    s_type                        StructureType
    p_next                        voidptr
    reduction_mode                SamplerReductionMode
} 

// PhysicalDeviceSamplerFilterMinmaxProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceSamplerFilterMinmaxProperties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    filter_minmax_single_component_formats Bool32
    filter_minmax_image_component_mapping Bool32
} 

// PhysicalDeviceVulkanMemoryModelFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceVulkanMemoryModelFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    vulkan_memory_model    Bool32
    vulkan_memory_model_device_scope Bool32
    vulkan_memory_model_availability_visibility_chains Bool32
} 

// PhysicalDeviceImagelessFramebufferFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceImagelessFramebufferFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    imageless_framebuffer  Bool32
} 

pub struct FramebufferAttachmentImageInfo {
mut:
    s_type                    StructureType
    p_next                    voidptr
    flags                     ImageCreateFlags
    usage                     ImageUsageFlags
    width                     u32
    height                    u32
    layer_count               u32
    view_format_count         u32
    p_view_formats            &Format
} 

// FramebufferAttachmentsCreateInfo extends VkFramebufferCreateInfo
pub struct FramebufferAttachmentsCreateInfo {
mut:
    s_type                                         StructureType
    p_next                                         voidptr
    attachment_image_info_count                    u32
    p_attachment_image_infos                       &FramebufferAttachmentImageInfo
} 

// RenderPassAttachmentBeginInfo extends VkRenderPassBeginInfo
pub struct RenderPassAttachmentBeginInfo {
mut:
    s_type                    StructureType
    p_next                    voidptr
    attachment_count          u32
    p_attachments             &C.ImageView
} 

// PhysicalDeviceUniformBufferStandardLayoutFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceUniformBufferStandardLayoutFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    uniform_buffer_standard_layout Bool32
} 

// PhysicalDeviceShaderSubgroupExtendedTypesFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderSubgroupExtendedTypesFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_subgroup_extended_types Bool32
} 

// PhysicalDeviceSeparateDepthStencilLayoutsFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceSeparateDepthStencilLayoutsFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    separate_depth_stencil_layouts Bool32
} 

// AttachmentReferenceStencilLayout extends VkAttachmentReference2
pub struct AttachmentReferenceStencilLayout {
mut:
    s_type                 StructureType
    p_next                 voidptr
    stencil_layout         ImageLayout
} 

// AttachmentDescriptionStencilLayout extends VkAttachmentDescription2
pub struct AttachmentDescriptionStencilLayout {
mut:
    s_type                 StructureType
    p_next                 voidptr
    stencil_initial_layout ImageLayout
    stencil_final_layout   ImageLayout
} 

// PhysicalDeviceHostQueryResetFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceHostQueryResetFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    host_query_reset       Bool32
} 

// PhysicalDeviceTimelineSemaphoreFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceTimelineSemaphoreFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    timeline_semaphore     Bool32
} 

// PhysicalDeviceTimelineSemaphoreProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceTimelineSemaphoreProperties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_timeline_semaphore_value_difference u64
} 

// SemaphoreTypeCreateInfo extends VkSemaphoreCreateInfo,VkPhysicalDeviceExternalSemaphoreInfo
pub struct SemaphoreTypeCreateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    semaphore_type         SemaphoreType
    initial_value          u64
} 

// TimelineSemaphoreSubmitInfo extends VkSubmitInfo,VkBindSparseInfo
pub struct TimelineSemaphoreSubmitInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    wait_semaphore_value_count u32
    p_wait_semaphore_values &u64
    signal_semaphore_value_count u32
    p_signal_semaphore_values &u64
} 

pub struct SemaphoreWaitInfo {
mut:
    s_type                      StructureType
    p_next                      voidptr
    flags                       SemaphoreWaitFlags
    semaphore_count             u32
    p_semaphores                &C.Semaphore
    p_values                    &u64
} 

pub struct SemaphoreSignalInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    semaphore              C.Semaphore
    value                  u64
} 

// PhysicalDeviceBufferDeviceAddressFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceBufferDeviceAddressFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    buffer_device_address  Bool32
    buffer_device_address_capture_replay Bool32
    buffer_device_address_multi_device Bool32
} 

pub struct BufferDeviceAddressInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    buffer                 C.Buffer
} 

// BufferOpaqueCaptureAddressCreateInfo extends VkBufferCreateInfo
pub struct BufferOpaqueCaptureAddressCreateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    opaque_capture_address u64
} 

// MemoryOpaqueCaptureAddressAllocateInfo extends VkMemoryAllocateInfo
pub struct MemoryOpaqueCaptureAddressAllocateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    opaque_capture_address u64
} 

pub struct DeviceMemoryOpaqueCaptureAddressInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    memory                 C.DeviceMemory
} 

type VkCmdDrawIndirectCount = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_indirect_count(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    count_buffer                                    C.Buffer,
    count_buffer_offset                             DeviceSize,
    max_draw_count                                  u32,
    stride                                          u32)  {
      f := VkCmdDrawIndirectCount((*loader_p).get_sym('vkCmdDrawIndirectCount'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawIndirectCount': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    count_buffer,
    count_buffer_offset,
    max_draw_count,
    stride)
}


type VkCmdDrawIndexedIndirectCount = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_indexed_indirect_count(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    count_buffer                                    C.Buffer,
    count_buffer_offset                             DeviceSize,
    max_draw_count                                  u32,
    stride                                          u32)  {
      f := VkCmdDrawIndexedIndirectCount((*loader_p).get_sym('vkCmdDrawIndexedIndirectCount'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawIndexedIndirectCount': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    count_buffer,
    count_buffer_offset,
    max_draw_count,
    stride)
}


type VkCreateRenderPass2 = fn (     C.Device,     &RenderPassCreateInfo2,     &AllocationCallbacks,     &C.RenderPass) Result

pub fn create_render_pass2(
    device                                          C.Device,
    p_create_info                                   &RenderPassCreateInfo2,
    p_allocator                                     &AllocationCallbacks,
    p_render_pass                                   &C.RenderPass) Result {
      f := VkCreateRenderPass2((*loader_p).get_sym('vkCreateRenderPass2'
    ) or { 
        println("Couldn't load symbol for 'vkCreateRenderPass2': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_render_pass)
}


type VkCmdBeginRenderPass2 = fn (     C.CommandBuffer,     &RenderPassBeginInfo,     &SubpassBeginInfo) 

pub fn cmd_begin_render_pass2(
    command_buffer                                  C.CommandBuffer,
    p_render_pass_begin                             &RenderPassBeginInfo,
    p_subpass_begin_info                            &SubpassBeginInfo)  {
      f := VkCmdBeginRenderPass2((*loader_p).get_sym('vkCmdBeginRenderPass2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBeginRenderPass2': ${err}")
        return 
    })
    f(
    command_buffer,
    p_render_pass_begin,
    p_subpass_begin_info)
}


type VkCmdNextSubpass2 = fn (     C.CommandBuffer,     &SubpassBeginInfo,     &SubpassEndInfo) 

pub fn cmd_next_subpass2(
    command_buffer                                  C.CommandBuffer,
    p_subpass_begin_info                            &SubpassBeginInfo,
    p_subpass_end_info                              &SubpassEndInfo)  {
      f := VkCmdNextSubpass2((*loader_p).get_sym('vkCmdNextSubpass2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdNextSubpass2': ${err}")
        return 
    })
    f(
    command_buffer,
    p_subpass_begin_info,
    p_subpass_end_info)
}


type VkCmdEndRenderPass2 = fn (     C.CommandBuffer,     &SubpassEndInfo) 

pub fn cmd_end_render_pass2(
    command_buffer                                  C.CommandBuffer,
    p_subpass_end_info                              &SubpassEndInfo)  {
      f := VkCmdEndRenderPass2((*loader_p).get_sym('vkCmdEndRenderPass2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEndRenderPass2': ${err}")
        return 
    })
    f(
    command_buffer,
    p_subpass_end_info)
}


type VkResetQueryPool = fn (     C.Device,     C.QueryPool,     u32,     u32) 

pub fn reset_query_pool(
    device                                          C.Device,
    query_pool                                      C.QueryPool,
    first_query                                     u32,
    query_count                                     u32)  {
      f := VkResetQueryPool((*loader_p).get_sym('vkResetQueryPool'
    ) or { 
        println("Couldn't load symbol for 'vkResetQueryPool': ${err}")
        return 
    })
    f(
    device,
    query_pool,
    first_query,
    query_count)
}


type VkGetSemaphoreCounterValue = fn (     C.Device,     C.Semaphore,     &u64) Result

pub fn get_semaphore_counter_value(
    device                                          C.Device,
    semaphore                                       C.Semaphore,
    p_value                                         &u64) Result {
      f := VkGetSemaphoreCounterValue((*loader_p).get_sym('vkGetSemaphoreCounterValue'
    ) or { 
        println("Couldn't load symbol for 'vkGetSemaphoreCounterValue': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    semaphore,
    p_value)
}


type VkWaitSemaphores = fn (     C.Device,     &SemaphoreWaitInfo,     u64) Result

pub fn wait_semaphores(
    device                                          C.Device,
    p_wait_info                                     &SemaphoreWaitInfo,
    timeout                                         u64) Result {
      f := VkWaitSemaphores((*loader_p).get_sym('vkWaitSemaphores'
    ) or { 
        println("Couldn't load symbol for 'vkWaitSemaphores': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_wait_info,
    timeout)
}


type VkSignalSemaphore = fn (     C.Device,     &SemaphoreSignalInfo) Result

pub fn signal_semaphore(
    device                                          C.Device,
    p_signal_info                                   &SemaphoreSignalInfo) Result {
      f := VkSignalSemaphore((*loader_p).get_sym('vkSignalSemaphore'
    ) or { 
        println("Couldn't load symbol for 'vkSignalSemaphore': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_signal_info)
}


type VkGetBufferDeviceAddress = fn (     C.Device,     &BufferDeviceAddressInfo) DeviceAddress

pub fn get_buffer_device_address(
    device                                          C.Device,
    p_info                                          &BufferDeviceAddressInfo) DeviceAddress {
      f := VkGetBufferDeviceAddress((*loader_p).get_sym("vkGetBufferDeviceAddress"
    ) or { 
        panic("Couldn't load symbol for 'vkGetBufferDeviceAddress': ${err}") })
    return f(
    device,
    p_info)
}


type VkGetBufferOpaqueCaptureAddress = fn (     C.Device,     &BufferDeviceAddressInfo) u64

pub fn get_buffer_opaque_capture_address(
    device                                          C.Device,
    p_info                                          &BufferDeviceAddressInfo) u64 {
      f := VkGetBufferOpaqueCaptureAddress((*loader_p).get_sym("vkGetBufferOpaqueCaptureAddress"
    ) or { 
        panic("Couldn't load symbol for 'vkGetBufferOpaqueCaptureAddress': ${err}") })
    return f(
    device,
    p_info)
}


type VkGetDeviceMemoryOpaqueCaptureAddress = fn (     C.Device,     &DeviceMemoryOpaqueCaptureAddressInfo) u64

pub fn get_device_memory_opaque_capture_address(
    device                                          C.Device,
    p_info                                          &DeviceMemoryOpaqueCaptureAddressInfo) u64 {
      f := VkGetDeviceMemoryOpaqueCaptureAddress((*loader_p).get_sym("vkGetDeviceMemoryOpaqueCaptureAddress"
    ) or { 
        panic("Couldn't load symbol for 'vkGetDeviceMemoryOpaqueCaptureAddress': ${err}") })
    return f(
    device,
    p_info)
}




// VK_VERSION_1_3 is a preprocessor guard. Do not pass it to API calls.
const version_1_3 = 1
// Vulkan 1.3 version number
pub const api_version_1_3 = make_api_version(0, 1, 3, 0)// Patch version should always be set to 0

pub type Flags64 = u64
pub type C.PrivateDataSlot = voidptr

pub enum PipelineCreationFeedbackFlagBits {
    pipeline_creation_feedback_valid_bit = int(0x00000001)
    pipeline_creation_feedback_application_pipeline_cache_hit_bit = int(0x00000002)
    pipeline_creation_feedback_base_pipeline_acceleration_bit = int(0x00000004)
    pipeline_creation_feedback_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type PipelineCreationFeedbackFlags = u32

pub enum ToolPurposeFlagBits {
    tool_purpose_validation_bit = int(0x00000001)
    tool_purpose_profiling_bit = int(0x00000002)
    tool_purpose_tracing_bit = int(0x00000004)
    tool_purpose_additional_features_bit = int(0x00000008)
    tool_purpose_modifying_features_bit = int(0x00000010)
    tool_purpose_debug_reporting_bit_ext = int(0x00000020)
    tool_purpose_debug_markers_bit_ext = int(0x00000040)
    tool_purpose_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type ToolPurposeFlags = u32
pub type PrivateDataSlotCreateFlags = u32
pub type PipelineStageFlags2 = u64

// Flag bits for PipelineStageFlagBits2
pub type PipelineStageFlagBits2 = u64
pub const pipeline_stage_2_none = u64(0)
pub const pipeline_stage_2_none_khr = pipeline_stage_2_none
pub const pipeline_stage_2_top_of_pipe_bit = u64(0x00000001)
pub const pipeline_stage_2_top_of_pipe_bit_khr = pipeline_stage_2_top_of_pipe_bit
pub const pipeline_stage_2_draw_indirect_bit = u64(0x00000002)
pub const pipeline_stage_2_draw_indirect_bit_khr = pipeline_stage_2_draw_indirect_bit
pub const pipeline_stage_2_vertex_input_bit = u64(0x00000004)
pub const pipeline_stage_2_vertex_input_bit_khr = u32(pipeline_stage_2_vertex_input_bit)
pub const pipeline_stage_2_vertex_shader_bit = u64(0x00000008)
pub const pipeline_stage_2_vertex_shader_bit_khr = pipeline_stage_2_vertex_shader_bit
pub const pipeline_stage_2_tessellation_control_shader_bit = u64(0x00000010)
pub const pipeline_stage_2_tessellation_control_shader_bit_khr = pipeline_stage_2_tessellation_control_shader_bit
pub const pipeline_stage_2_tessellation_evaluation_shader_bit = u64(0x00000020)
pub const pipeline_stage_2_tessellation_evaluation_shader_bit_khr = u32(pipeline_stage_2_tessellation_evaluation_shader_bit)
pub const pipeline_stage_2_geometry_shader_bit = u64(0x00000040)
pub const pipeline_stage_2_geometry_shader_bit_khr = pipeline_stage_2_geometry_shader_bit
pub const pipeline_stage_2_fragment_shader_bit = u64(0x00000080)
pub const pipeline_stage_2_fragment_shader_bit_khr = pipeline_stage_2_fragment_shader_bit
pub const pipeline_stage_2_early_fragment_tests_bit = u64(0x00000100)
pub const pipeline_stage_2_early_fragment_tests_bit_khr = pipeline_stage_2_early_fragment_tests_bit
pub const pipeline_stage_2_late_fragment_tests_bit = u64(0x00000200)
pub const pipeline_stage_2_late_fragment_tests_bit_khr = pipeline_stage_2_late_fragment_tests_bit
pub const pipeline_stage_2_color_attachment_output_bit = u64(0x00000400)
pub const pipeline_stage_2_color_attachment_output_bit_khr = u32(pipeline_stage_2_color_attachment_output_bit)
pub const pipeline_stage_2_compute_shader_bit = u64(0x00000800)
pub const pipeline_stage_2_compute_shader_bit_khr = u32(pipeline_stage_2_compute_shader_bit)
pub const pipeline_stage_2_all_transfer_bit = u64(0x00001000)
pub const pipeline_stage_2_all_transfer_bit_khr = pipeline_stage_2_all_transfer_bit
pub const pipeline_stage_2_transfer_bit = pipeline_stage_2_all_transfer_bit_khr
pub const pipeline_stage_2_transfer_bit_khr = pipeline_stage_2_all_transfer_bit
pub const pipeline_stage_2_bottom_of_pipe_bit = u64(0x00002000)
pub const pipeline_stage_2_bottom_of_pipe_bit_khr = pipeline_stage_2_bottom_of_pipe_bit
pub const pipeline_stage_2_host_bit = u64(0x00004000)
pub const pipeline_stage_2_host_bit_khr = pipeline_stage_2_host_bit
pub const pipeline_stage_2_all_graphics_bit = u64(0x00008000)
pub const pipeline_stage_2_all_graphics_bit_khr = pipeline_stage_2_all_graphics_bit
pub const pipeline_stage_2_all_commands_bit = u64(0x00010000)
pub const pipeline_stage_2_all_commands_bit_khr = pipeline_stage_2_all_commands_bit
pub const pipeline_stage_2_copy_bit = u64(0x100000000)
pub const pipeline_stage_2_copy_bit_khr = pipeline_stage_2_copy_bit
pub const pipeline_stage_2_resolve_bit = u64(0x200000000)
pub const pipeline_stage_2_resolve_bit_khr = pipeline_stage_2_resolve_bit
pub const pipeline_stage_2_blit_bit = u64(0x400000000)
pub const pipeline_stage_2_blit_bit_khr = pipeline_stage_2_blit_bit
pub const pipeline_stage_2_clear_bit = u64(0x800000000)
pub const pipeline_stage_2_clear_bit_khr = pipeline_stage_2_clear_bit
pub const pipeline_stage_2_index_input_bit = u64(0x1000000000)
pub const pipeline_stage_2_index_input_bit_khr = u32(pipeline_stage_2_index_input_bit)
pub const pipeline_stage_2_vertex_attribute_input_bit = u64(0x2000000000)
pub const pipeline_stage_2_vertex_attribute_input_bit_khr = u32(pipeline_stage_2_vertex_attribute_input_bit)
pub const pipeline_stage_2_pre_rasterization_shaders_bit = u64(0x4000000000)
pub const pipeline_stage_2_pre_rasterization_shaders_bit_khr = pipeline_stage_2_pre_rasterization_shaders_bit
pub const pipeline_stage_2_video_decode_bit_khr = u64(0x04000000)
pub const pipeline_stage_2_transform_feedback_bit_ext = u64(0x01000000)
pub const pipeline_stage_2_conditional_rendering_bit_ext = u64(0x00040000)
pub const pipeline_stage_2_command_preprocess_bit_nv = u64(0x00020000)
pub const pipeline_stage_2_fragment_shading_rate_attachment_bit_khr = u64(0x00400000)
pub const pipeline_stage_2_shading_rate_image_bit_nv = pipeline_stage_2_fragment_shading_rate_attachment_bit_khr
pub const pipeline_stage_2_acceleration_structure_build_bit_khr = u64(0x02000000)
pub const pipeline_stage_2_ray_tracing_shader_bit_khr = u64(0x00200000)
pub const pipeline_stage_2_ray_tracing_shader_bit_nv = pipeline_stage_2_ray_tracing_shader_bit_khr
pub const pipeline_stage_2_acceleration_structure_build_bit_nv = u32(pipeline_stage_2_acceleration_structure_build_bit_khr)
pub const pipeline_stage_2_fragment_density_process_bit_ext = u64(0x00800000)
pub const pipeline_stage_2_task_shader_bit_nv = pipeline_stage_2_task_shader_bit_ext
pub const pipeline_stage_2_mesh_shader_bit_nv = pipeline_stage_2_mesh_shader_bit_ext
pub const pipeline_stage_2_task_shader_bit_ext = u64(0x00080000)
pub const pipeline_stage_2_mesh_shader_bit_ext = u64(0x00100000)
pub const pipeline_stage_2_subpass_shader_bit_huawei = u64(0x8000000000)
pub const pipeline_stage_2_subpass_shading_bit_huawei = u32(pipeline_stage_2_subpass_shader_bit_huawei)
pub const pipeline_stage_2_invocation_mask_bit_huawei = u64(0x10000000000)
pub const pipeline_stage_2_acceleration_structure_copy_bit_khr = u64(0x10000000)
pub const pipeline_stage_2_micromap_build_bit_ext = u64(0x40000000)
pub const pipeline_stage_2_cluster_culling_shader_bit_huawei = u64(0x20000000000)
pub const pipeline_stage_2_optical_flow_bit_nv = u64(0x20000000)


pub type AccessFlags2 = u64

// Flag bits for AccessFlagBits2
pub type AccessFlagBits2 = u64
pub const access_2_none = u64(0)
pub const access_2_none_khr = access_2_none
pub const access_2_indirect_command_read_bit = u64(0x00000001)
pub const access_2_indirect_command_read_bit_khr = access_2_indirect_command_read_bit
pub const access_2_index_read_bit = u64(0x00000002)
pub const access_2_index_read_bit_khr = access_2_index_read_bit
pub const access_2_vertex_attribute_read_bit = u64(0x00000004)
pub const access_2_vertex_attribute_read_bit_khr = u32(access_2_vertex_attribute_read_bit)
pub const access_2_uniform_read_bit = u64(0x00000008)
pub const access_2_uniform_read_bit_khr = u32(access_2_uniform_read_bit)
pub const access_2_input_attachment_read_bit = u64(0x00000010)
pub const access_2_input_attachment_read_bit_khr = u32(access_2_input_attachment_read_bit)
pub const access_2_shader_read_bit = u64(0x00000020)
pub const access_2_shader_read_bit_khr = access_2_shader_read_bit
pub const access_2_shader_write_bit = u64(0x00000040)
pub const access_2_shader_write_bit_khr = access_2_shader_write_bit
pub const access_2_color_attachment_read_bit = u64(0x00000080)
pub const access_2_color_attachment_read_bit_khr = access_2_color_attachment_read_bit
pub const access_2_color_attachment_write_bit = u64(0x00000100)
pub const access_2_color_attachment_write_bit_khr = access_2_color_attachment_write_bit
pub const access_2_depth_stencil_attachment_read_bit = u64(0x00000200)
pub const access_2_depth_stencil_attachment_read_bit_khr = access_2_depth_stencil_attachment_read_bit
pub const access_2_depth_stencil_attachment_write_bit = u64(0x00000400)
pub const access_2_depth_stencil_attachment_write_bit_khr = access_2_depth_stencil_attachment_write_bit
pub const access_2_transfer_read_bit = u64(0x00000800)
pub const access_2_transfer_read_bit_khr = access_2_transfer_read_bit
pub const access_2_transfer_write_bit = u64(0x00001000)
pub const access_2_transfer_write_bit_khr = access_2_transfer_write_bit
pub const access_2_host_read_bit = u64(0x00002000)
pub const access_2_host_read_bit_khr = access_2_host_read_bit
pub const access_2_host_write_bit = u64(0x00004000)
pub const access_2_host_write_bit_khr = access_2_host_write_bit
pub const access_2_memory_read_bit = u64(0x00008000)
pub const access_2_memory_read_bit_khr = access_2_memory_read_bit
pub const access_2_memory_write_bit = u64(0x00010000)
pub const access_2_memory_write_bit_khr = access_2_memory_write_bit
pub const access_2_shader_sampled_read_bit = u64(0x100000000)
pub const access_2_shader_sampled_read_bit_khr = access_2_shader_sampled_read_bit
pub const access_2_shader_storage_read_bit = u64(0x200000000)
pub const access_2_shader_storage_read_bit_khr = access_2_shader_storage_read_bit
pub const access_2_shader_storage_write_bit = u64(0x400000000)
pub const access_2_shader_storage_write_bit_khr = access_2_shader_storage_write_bit
pub const access_2_video_decode_read_bit_khr = u64(0x800000000)
pub const access_2_video_decode_write_bit_khr = u64(0x1000000000)
pub const access_2_transform_feedback_write_bit_ext = u64(0x02000000)
pub const access_2_transform_feedback_counter_read_bit_ext = u64(0x04000000)
pub const access_2_transform_feedback_counter_write_bit_ext = u64(0x08000000)
pub const access_2_conditional_rendering_read_bit_ext = u64(0x00100000)
pub const access_2_command_preprocess_read_bit_nv = u64(0x00020000)
pub const access_2_command_preprocess_write_bit_nv = u64(0x00040000)
pub const access_2_fragment_shading_rate_attachment_read_bit_khr = u64(0x00800000)
pub const access_2_shading_rate_image_read_bit_nv = access_2_fragment_shading_rate_attachment_read_bit_khr
pub const access_2_acceleration_structure_read_bit_khr = u64(0x00200000)
pub const access_2_acceleration_structure_write_bit_khr = u64(0x00400000)
pub const access_2_acceleration_structure_read_bit_nv = u32(access_2_acceleration_structure_read_bit_khr)
pub const access_2_acceleration_structure_write_bit_nv = u32(access_2_acceleration_structure_write_bit_khr)
pub const access_2_fragment_density_map_read_bit_ext = u64(0x01000000)
pub const access_2_color_attachment_read_noncoherent_bit_ext = u64(0x00080000)
pub const access_2_descriptor_buffer_read_bit_ext = u64(0x20000000000)
pub const access_2_invocation_mask_read_bit_huawei = u64(0x8000000000)
pub const access_2_shader_binding_table_read_bit_khr = u64(0x10000000000)
pub const access_2_micromap_read_bit_ext = u64(0x100000000000)
pub const access_2_micromap_write_bit_ext = u64(0x200000000000)
pub const access_2_optical_flow_read_bit_nv = u64(0x40000000000)
pub const access_2_optical_flow_write_bit_nv = u64(0x80000000000)



pub enum SubmitFlagBits {
    submit_protected_bit = int(0x00000001)
    submit_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type SubmitFlags = u32

pub enum RenderingFlagBits {
    rendering_contents_secondary_command_buffers_bit = int(0x00000001)
    rendering_suspending_bit = int(0x00000002)
    rendering_resuming_bit = int(0x00000004)
    rendering_contents_inline_bit_ext = int(0x00000010)
    rendering_enable_legacy_dithering_bit_ext = int(0x00000008)
    rendering_flag_bits_max_enum = int(0x7FFFFFFF)
}

pub type RenderingFlags = u32
pub type FormatFeatureFlags2 = u64

// Flag bits for FormatFeatureFlagBits2
pub type FormatFeatureFlagBits2 = u64
pub const format_feature_2_sampled_image_bit = u64(0x00000001)
pub const format_feature_2_sampled_image_bit_khr = u32(format_feature_2_sampled_image_bit)
pub const format_feature_2_storage_image_bit = u64(0x00000002)
pub const format_feature_2_storage_image_bit_khr = u32(format_feature_2_storage_image_bit)
pub const format_feature_2_storage_image_atomic_bit = u64(0x00000004)
pub const format_feature_2_storage_image_atomic_bit_khr = u32(format_feature_2_storage_image_atomic_bit)
pub const format_feature_2_uniform_texel_buffer_bit = u64(0x00000008)
pub const format_feature_2_uniform_texel_buffer_bit_khr = u32(format_feature_2_uniform_texel_buffer_bit)
pub const format_feature_2_storage_texel_buffer_bit = u64(0x00000010)
pub const format_feature_2_storage_texel_buffer_bit_khr = u32(format_feature_2_storage_texel_buffer_bit)
pub const format_feature_2_storage_texel_buffer_atomic_bit = u64(0x00000020)
pub const format_feature_2_storage_texel_buffer_atomic_bit_khr = u32(format_feature_2_storage_texel_buffer_atomic_bit)
pub const format_feature_2_vertex_buffer_bit = u64(0x00000040)
pub const format_feature_2_vertex_buffer_bit_khr = u32(format_feature_2_vertex_buffer_bit)
pub const format_feature_2_color_attachment_bit = u64(0x00000080)
pub const format_feature_2_color_attachment_bit_khr = u32(format_feature_2_color_attachment_bit)
pub const format_feature_2_color_attachment_blend_bit = u64(0x00000100)
pub const format_feature_2_color_attachment_blend_bit_khr = u32(format_feature_2_color_attachment_blend_bit)
pub const format_feature_2_depth_stencil_attachment_bit = u64(0x00000200)
pub const format_feature_2_depth_stencil_attachment_bit_khr = u32(format_feature_2_depth_stencil_attachment_bit)
pub const format_feature_2_blit_src_bit = u64(0x00000400)
pub const format_feature_2_blit_src_bit_khr = u32(format_feature_2_blit_src_bit)
pub const format_feature_2_blit_dst_bit = u64(0x00000800)
pub const format_feature_2_blit_dst_bit_khr = u32(format_feature_2_blit_dst_bit)
pub const format_feature_2_sampled_image_filter_linear_bit = u64(0x00001000)
pub const format_feature_2_sampled_image_filter_linear_bit_khr = u32(format_feature_2_sampled_image_filter_linear_bit)
pub const format_feature_2_sampled_image_filter_cubic_bit = u64(0x00002000)
pub const format_feature_2_sampled_image_filter_cubic_bit_ext = u32(format_feature_2_sampled_image_filter_cubic_bit)
pub const format_feature_2_transfer_src_bit = u64(0x00004000)
pub const format_feature_2_transfer_src_bit_khr = u32(format_feature_2_transfer_src_bit)
pub const format_feature_2_transfer_dst_bit = u64(0x00008000)
pub const format_feature_2_transfer_dst_bit_khr = u32(format_feature_2_transfer_dst_bit)
pub const format_feature_2_sampled_image_filter_minmax_bit = u64(0x00010000)
pub const format_feature_2_sampled_image_filter_minmax_bit_khr = u32(format_feature_2_sampled_image_filter_minmax_bit)
pub const format_feature_2_midpoint_chroma_samples_bit = u64(0x00020000)
pub const format_feature_2_midpoint_chroma_samples_bit_khr = u32(format_feature_2_midpoint_chroma_samples_bit)
pub const format_feature_2_sampled_image_ycbcr_conversion_linear_filter_bit = u64(0x00040000)
pub const format_feature_2_sampled_image_ycbcr_conversion_linear_filter_bit_khr = u32(format_feature_2_sampled_image_ycbcr_conversion_linear_filter_bit)
pub const format_feature_2_sampled_image_ycbcr_conversion_separate_reconstruction_filter_bit = u64(0x00080000)
pub const format_feature_2_sampled_image_ycbcr_conversion_separate_reconstruction_filter_bit_khr = u32(format_feature_2_sampled_image_ycbcr_conversion_separate_reconstruction_filter_bit)
pub const format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_bit = u64(0x00100000)
pub const format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_bit_khr = u32(format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_bit)
pub const format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_forceable_bit = u64(0x00200000)
pub const format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_forceable_bit_khr = u32(format_feature_2_sampled_image_ycbcr_conversion_chroma_reconstruction_explicit_forceable_bit)
pub const format_feature_2_disjoint_bit = u64(0x00400000)
pub const format_feature_2_disjoint_bit_khr = u32(format_feature_2_disjoint_bit)
pub const format_feature_2_cosited_chroma_samples_bit = u64(0x00800000)
pub const format_feature_2_cosited_chroma_samples_bit_khr = u32(format_feature_2_cosited_chroma_samples_bit)
pub const format_feature_2_storage_read_without_format_bit = u64(0x80000000)
pub const format_feature_2_storage_read_without_format_bit_khr = u32(format_feature_2_storage_read_without_format_bit)
pub const format_feature_2_storage_write_without_format_bit = u64(0x100000000)
pub const format_feature_2_storage_write_without_format_bit_khr = u32(format_feature_2_storage_write_without_format_bit)
pub const format_feature_2_sampled_image_depth_comparison_bit = u64(0x200000000)
pub const format_feature_2_sampled_image_depth_comparison_bit_khr = u32(format_feature_2_sampled_image_depth_comparison_bit)
pub const format_feature_2_video_decode_output_bit_khr = u64(0x02000000)
pub const format_feature_2_video_decode_dpb_bit_khr = u64(0x04000000)
pub const format_feature_2_acceleration_structure_vertex_buffer_bit_khr = u64(0x20000000)
pub const format_feature_2_fragment_density_map_bit_ext = u64(0x01000000)
pub const format_feature_2_fragment_shading_rate_attachment_bit_khr = u64(0x40000000)
pub const format_feature_2_host_image_transfer_bit_ext = u64(0x400000000000)
pub const format_feature_2_linear_color_attachment_bit_nv = u64(0x4000000000)
pub const format_feature_2_weight_image_bit_qcom = u64(0x400000000)
pub const format_feature_2_weight_sampled_image_bit_qcom = u64(0x800000000)
pub const format_feature_2_block_matching_bit_qcom = u64(0x1000000000)
pub const format_feature_2_box_filter_sampled_bit_qcom = u64(0x2000000000)
pub const format_feature_2_optical_flow_image_bit_nv = u64(0x10000000000)
pub const format_feature_2_optical_flow_vector_bit_nv = u64(0x20000000000)
pub const format_feature_2_optical_flow_cost_bit_nv = u64(0x40000000000)


// PhysicalDeviceVulkan13Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceVulkan13Features {
mut:
    s_type                 StructureType
    p_next                 voidptr
    robust_image_access    Bool32
    inline_uniform_block   Bool32
    descriptor_binding_inline_uniform_block_update_after_bind Bool32
    pipeline_creation_cache_control Bool32
    private_data           Bool32
    shader_demote_to_helper_invocation Bool32
    shader_terminate_invocation Bool32
    subgroup_size_control  Bool32
    compute_full_subgroups Bool32
    synchronization2       Bool32
    texture_compression_astc_hdr Bool32
    shader_zero_initialize_workgroup_memory Bool32
    dynamic_rendering      Bool32
    shader_integer_dot_product Bool32
    maintenance4           Bool32
} 

// PhysicalDeviceVulkan13Properties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceVulkan13Properties {
mut:
    s_type                    StructureType
    p_next                    voidptr
    min_subgroup_size         u32
    max_subgroup_size         u32
    max_compute_workgroup_subgroups u32
    required_subgroup_size_stages ShaderStageFlags
    max_inline_uniform_block_size u32
    max_per_stage_descriptor_inline_uniform_blocks u32
    max_per_stage_descriptor_update_after_bind_inline_uniform_blocks u32
    max_descriptor_set_inline_uniform_blocks u32
    max_descriptor_set_update_after_bind_inline_uniform_blocks u32
    max_inline_uniform_total_size u32
    integer_dot_product8_bit_unsigned_accelerated Bool32
    integer_dot_product8_bit_signed_accelerated Bool32
    integer_dot_product8_bit_mixed_signedness_accelerated Bool32
    integer_dot_product4x8_bit_packed_unsigned_accelerated Bool32
    integer_dot_product4x8_bit_packed_signed_accelerated Bool32
    integer_dot_product4x8_bit_packed_mixed_signedness_accelerated Bool32
    integer_dot_product16_bit_unsigned_accelerated Bool32
    integer_dot_product16_bit_signed_accelerated Bool32
    integer_dot_product16_bit_mixed_signedness_accelerated Bool32
    integer_dot_product32_bit_unsigned_accelerated Bool32
    integer_dot_product32_bit_signed_accelerated Bool32
    integer_dot_product32_bit_mixed_signedness_accelerated Bool32
    integer_dot_product64_bit_unsigned_accelerated Bool32
    integer_dot_product64_bit_signed_accelerated Bool32
    integer_dot_product64_bit_mixed_signedness_accelerated Bool32
    integer_dot_product_accumulating_saturating8_bit_unsigned_accelerated Bool32
    integer_dot_product_accumulating_saturating8_bit_signed_accelerated Bool32
    integer_dot_product_accumulating_saturating8_bit_mixed_signedness_accelerated Bool32
    integer_dot_product_accumulating_saturating4x8_bit_packed_unsigned_accelerated Bool32
    integer_dot_product_accumulating_saturating4x8_bit_packed_signed_accelerated Bool32
    integer_dot_product_accumulating_saturating4x8_bit_packed_mixed_signedness_accelerated Bool32
    integer_dot_product_accumulating_saturating16_bit_unsigned_accelerated Bool32
    integer_dot_product_accumulating_saturating16_bit_signed_accelerated Bool32
    integer_dot_product_accumulating_saturating16_bit_mixed_signedness_accelerated Bool32
    integer_dot_product_accumulating_saturating32_bit_unsigned_accelerated Bool32
    integer_dot_product_accumulating_saturating32_bit_signed_accelerated Bool32
    integer_dot_product_accumulating_saturating32_bit_mixed_signedness_accelerated Bool32
    integer_dot_product_accumulating_saturating64_bit_unsigned_accelerated Bool32
    integer_dot_product_accumulating_saturating64_bit_signed_accelerated Bool32
    integer_dot_product_accumulating_saturating64_bit_mixed_signedness_accelerated Bool32
    storage_texel_buffer_offset_alignment_bytes DeviceSize
    storage_texel_buffer_offset_single_texel_alignment Bool32
    uniform_texel_buffer_offset_alignment_bytes DeviceSize
    uniform_texel_buffer_offset_single_texel_alignment Bool32
    max_buffer_size           DeviceSize
} 

pub struct PipelineCreationFeedback {
mut:
    flags                                  PipelineCreationFeedbackFlags
    duration                               u64
} 

// PipelineCreationFeedbackCreateInfo extends VkGraphicsPipelineCreateInfo,VkComputePipelineCreateInfo,VkRayTracingPipelineCreateInfoNV,VkRayTracingPipelineCreateInfoKHR,VkExecutionGraphPipelineCreateInfoAMDX
pub struct PipelineCreationFeedbackCreateInfo {
mut:
    s_type                             StructureType
    p_next                             voidptr
    p_pipeline_creation_feedback       &PipelineCreationFeedback
    pipeline_stage_creation_feedback_count u32
    p_pipeline_stage_creation_feedbacks &PipelineCreationFeedback
} 

// PhysicalDeviceShaderTerminateInvocationFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderTerminateInvocationFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_terminate_invocation Bool32
} 

pub struct PhysicalDeviceToolProperties {
mut:
    s_type                    StructureType
    p_next                    voidptr
    name                      []char
    version                   []char
    purposes                  ToolPurposeFlags
    description               []char
    layer                     []char
} 

// PhysicalDeviceShaderDemoteToHelperInvocationFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderDemoteToHelperInvocationFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_demote_to_helper_invocation Bool32
} 

// PhysicalDevicePrivateDataFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePrivateDataFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    private_data           Bool32
} 

// DevicePrivateDataCreateInfo extends VkDeviceCreateInfo
pub struct DevicePrivateDataCreateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    private_data_slot_request_count u32
} 

pub struct PrivateDataSlotCreateInfo {
mut:
    s_type                              StructureType
    p_next                              voidptr
    flags                               PrivateDataSlotCreateFlags
} 

// PhysicalDevicePipelineCreationCacheControlFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePipelineCreationCacheControlFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pipeline_creation_cache_control Bool32
} 

// MemoryBarrier2 extends VkSubpassDependency2
pub struct MemoryBarrier2 {
mut:
    s_type                       StructureType
    p_next                       voidptr
    src_stage_mask               PipelineStageFlags2
    src_access_mask              AccessFlags2
    dst_stage_mask               PipelineStageFlags2
    dst_access_mask              AccessFlags2
} 

pub struct BufferMemoryBarrier2 {
mut:
    s_type                       StructureType
    p_next                       voidptr
    src_stage_mask               PipelineStageFlags2
    src_access_mask              AccessFlags2
    dst_stage_mask               PipelineStageFlags2
    dst_access_mask              AccessFlags2
    src_queue_family_index       u32
    dst_queue_family_index       u32
    buffer                       C.Buffer
    offset                       DeviceSize
    size                         DeviceSize
} 

pub struct ImageMemoryBarrier2 {
mut:
    s_type                         StructureType
    p_next                         voidptr
    src_stage_mask                 PipelineStageFlags2
    src_access_mask                AccessFlags2
    dst_stage_mask                 PipelineStageFlags2
    dst_access_mask                AccessFlags2
    old_layout                     ImageLayout
    new_layout                     ImageLayout
    src_queue_family_index         u32
    dst_queue_family_index         u32
    image                          C.Image
    subresource_range              ImageSubresourceRange
} 

pub struct DependencyInfo {
mut:
    s_type                               StructureType
    p_next                               voidptr
    dependency_flags                     DependencyFlags
    memory_barrier_count                 u32
    p_memory_barriers                    &MemoryBarrier2
    buffer_memory_barrier_count          u32
    p_buffer_memory_barriers             &BufferMemoryBarrier2
    image_memory_barrier_count           u32
    p_image_memory_barriers              &ImageMemoryBarrier2
} 

pub struct SemaphoreSubmitInfo {
mut:
    s_type                       StructureType
    p_next                       voidptr
    semaphore                    C.Semaphore
    value                        u64
    stage_mask                   PipelineStageFlags2
    device_index                 u32
} 

pub struct CommandBufferSubmitInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    command_buffer         C.CommandBuffer
    device_mask            u32
} 

pub struct SubmitInfo2 {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    flags                                   SubmitFlags
    wait_semaphore_info_count               u32
    p_wait_semaphore_infos                  &SemaphoreSubmitInfo
    command_buffer_info_count               u32
    p_command_buffer_infos                  &CommandBufferSubmitInfo
    signal_semaphore_info_count             u32
    p_signal_semaphore_infos                &SemaphoreSubmitInfo
} 

// PhysicalDeviceSynchronization2Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceSynchronization2Features {
mut:
    s_type                 StructureType
    p_next                 voidptr
    synchronization2       Bool32
} 

// PhysicalDeviceZeroInitializeWorkgroupMemoryFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceZeroInitializeWorkgroupMemoryFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_zero_initialize_workgroup_memory Bool32
} 

// PhysicalDeviceImageRobustnessFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceImageRobustnessFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    robust_image_access    Bool32
} 

pub struct BufferCopy2 {
mut:
    s_type                 StructureType
    p_next                 voidptr
    src_offset             DeviceSize
    dst_offset             DeviceSize
    size                   DeviceSize
} 

pub struct CopyBufferInfo2 {
mut:
    s_type                      StructureType
    p_next                      voidptr
    src_buffer                  C.Buffer
    dst_buffer                  C.Buffer
    region_count                u32
    p_regions                   &BufferCopy2
} 

pub struct ImageCopy2 {
mut:
    s_type                          StructureType
    p_next                          voidptr
    src_subresource                 ImageSubresourceLayers
    src_offset                      Offset3D
    dst_subresource                 ImageSubresourceLayers
    dst_offset                      Offset3D
    extent                          Extent3D
} 

pub struct CopyImageInfo2 {
mut:
    s_type                     StructureType
    p_next                     voidptr
    src_image                  C.Image
    src_image_layout           ImageLayout
    dst_image                  C.Image
    dst_image_layout           ImageLayout
    region_count               u32
    p_regions                  &ImageCopy2
} 

pub struct BufferImageCopy2 {
mut:
    s_type                          StructureType
    p_next                          voidptr
    buffer_offset                   DeviceSize
    buffer_row_length               u32
    buffer_image_height             u32
    image_subresource               ImageSubresourceLayers
    image_offset                    Offset3D
    image_extent                    Extent3D
} 

pub struct CopyBufferToImageInfo2 {
mut:
    s_type                           StructureType
    p_next                           voidptr
    src_buffer                       C.Buffer
    dst_image                        C.Image
    dst_image_layout                 ImageLayout
    region_count                     u32
    p_regions                        &BufferImageCopy2
} 

pub struct CopyImageToBufferInfo2 {
mut:
    s_type                           StructureType
    p_next                           voidptr
    src_image                        C.Image
    src_image_layout                 ImageLayout
    dst_buffer                       C.Buffer
    region_count                     u32
    p_regions                        &BufferImageCopy2
} 

pub struct ImageBlit2 {
mut:
    s_type                          StructureType
    p_next                          voidptr
    src_subresource                 ImageSubresourceLayers
    src_offsets                     []Offset3D
    dst_subresource                 ImageSubresourceLayers
    dst_offsets                     []Offset3D
} 

pub struct BlitImageInfo2 {
mut:
    s_type                     StructureType
    p_next                     voidptr
    src_image                  C.Image
    src_image_layout           ImageLayout
    dst_image                  C.Image
    dst_image_layout           ImageLayout
    region_count               u32
    p_regions                  &ImageBlit2
    filter                     Filter
} 

pub struct ImageResolve2 {
mut:
    s_type                          StructureType
    p_next                          voidptr
    src_subresource                 ImageSubresourceLayers
    src_offset                      Offset3D
    dst_subresource                 ImageSubresourceLayers
    dst_offset                      Offset3D
    extent                          Extent3D
} 

pub struct ResolveImageInfo2 {
mut:
    s_type                        StructureType
    p_next                        voidptr
    src_image                     C.Image
    src_image_layout              ImageLayout
    dst_image                     C.Image
    dst_image_layout              ImageLayout
    region_count                  u32
    p_regions                     &ImageResolve2
} 

// PhysicalDeviceSubgroupSizeControlFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceSubgroupSizeControlFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    subgroup_size_control  Bool32
    compute_full_subgroups Bool32
} 

// PhysicalDeviceSubgroupSizeControlProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceSubgroupSizeControlProperties {
mut:
    s_type                    StructureType
    p_next                    voidptr
    min_subgroup_size         u32
    max_subgroup_size         u32
    max_compute_workgroup_subgroups u32
    required_subgroup_size_stages ShaderStageFlags
} 

// PipelineShaderStageRequiredSubgroupSizeCreateInfo extends VkPipelineShaderStageCreateInfo,VkShaderCreateInfoEXT
pub struct PipelineShaderStageRequiredSubgroupSizeCreateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    required_subgroup_size u32
} 

// PhysicalDeviceInlineUniformBlockFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceInlineUniformBlockFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    inline_uniform_block   Bool32
    descriptor_binding_inline_uniform_block_update_after_bind Bool32
} 

// PhysicalDeviceInlineUniformBlockProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceInlineUniformBlockProperties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_inline_uniform_block_size u32
    max_per_stage_descriptor_inline_uniform_blocks u32
    max_per_stage_descriptor_update_after_bind_inline_uniform_blocks u32
    max_descriptor_set_inline_uniform_blocks u32
    max_descriptor_set_update_after_bind_inline_uniform_blocks u32
} 

// WriteDescriptorSetInlineUniformBlock extends VkWriteDescriptorSet
pub struct WriteDescriptorSetInlineUniformBlock {
mut:
    s_type                 StructureType
    p_next                 voidptr
    data_size              u32
    p_data                 voidptr
} 

// DescriptorPoolInlineUniformBlockCreateInfo extends VkDescriptorPoolCreateInfo
pub struct DescriptorPoolInlineUniformBlockCreateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_inline_uniform_block_bindings u32
} 

// PhysicalDeviceTextureCompressionASTCHDRFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceTextureCompressionASTCHDRFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    texture_compression_astc_hdr Bool32
} 

pub struct RenderingAttachmentInfo {
mut:
    s_type                       StructureType
    p_next                       voidptr
    image_view                   C.ImageView
    image_layout                 ImageLayout
    resolve_mode                 ResolveModeFlagBits
    resolve_image_view           C.ImageView
    resolve_image_layout         ImageLayout
    load_op                      AttachmentLoadOp
    store_op                     AttachmentStoreOp
    clear_value                  ClearValue
} 

pub struct RenderingInfo {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    flags                                   RenderingFlags
    render_area                             Rect2D
    layer_count                             u32
    view_mask                               u32
    color_attachment_count                  u32
    p_color_attachments                     &RenderingAttachmentInfo
    p_depth_attachment                      &RenderingAttachmentInfo
    p_stencil_attachment                    &RenderingAttachmentInfo
} 

// PipelineRenderingCreateInfo extends VkGraphicsPipelineCreateInfo
pub struct PipelineRenderingCreateInfo {
mut:
    s_type                 StructureType
    p_next                 voidptr
    view_mask              u32
    color_attachment_count u32
    p_color_attachment_formats &Format
    depth_attachment_format Format
    stencil_attachment_format Format
} 

// PhysicalDeviceDynamicRenderingFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDynamicRenderingFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    dynamic_rendering      Bool32
} 

// CommandBufferInheritanceRenderingInfo extends VkCommandBufferInheritanceInfo
pub struct CommandBufferInheritanceRenderingInfo {
mut:
    s_type                       StructureType
    p_next                       voidptr
    flags                        RenderingFlags
    view_mask                    u32
    color_attachment_count       u32
    p_color_attachment_formats   &Format
    depth_attachment_format      Format
    stencil_attachment_format    Format
    rasterization_samples        SampleCountFlagBits
} 

// PhysicalDeviceShaderIntegerDotProductFeatures extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderIntegerDotProductFeatures {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_integer_dot_product Bool32
} 

// PhysicalDeviceShaderIntegerDotProductProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceShaderIntegerDotProductProperties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    integer_dot_product8_bit_unsigned_accelerated Bool32
    integer_dot_product8_bit_signed_accelerated Bool32
    integer_dot_product8_bit_mixed_signedness_accelerated Bool32
    integer_dot_product4x8_bit_packed_unsigned_accelerated Bool32
    integer_dot_product4x8_bit_packed_signed_accelerated Bool32
    integer_dot_product4x8_bit_packed_mixed_signedness_accelerated Bool32
    integer_dot_product16_bit_unsigned_accelerated Bool32
    integer_dot_product16_bit_signed_accelerated Bool32
    integer_dot_product16_bit_mixed_signedness_accelerated Bool32
    integer_dot_product32_bit_unsigned_accelerated Bool32
    integer_dot_product32_bit_signed_accelerated Bool32
    integer_dot_product32_bit_mixed_signedness_accelerated Bool32
    integer_dot_product64_bit_unsigned_accelerated Bool32
    integer_dot_product64_bit_signed_accelerated Bool32
    integer_dot_product64_bit_mixed_signedness_accelerated Bool32
    integer_dot_product_accumulating_saturating8_bit_unsigned_accelerated Bool32
    integer_dot_product_accumulating_saturating8_bit_signed_accelerated Bool32
    integer_dot_product_accumulating_saturating8_bit_mixed_signedness_accelerated Bool32
    integer_dot_product_accumulating_saturating4x8_bit_packed_unsigned_accelerated Bool32
    integer_dot_product_accumulating_saturating4x8_bit_packed_signed_accelerated Bool32
    integer_dot_product_accumulating_saturating4x8_bit_packed_mixed_signedness_accelerated Bool32
    integer_dot_product_accumulating_saturating16_bit_unsigned_accelerated Bool32
    integer_dot_product_accumulating_saturating16_bit_signed_accelerated Bool32
    integer_dot_product_accumulating_saturating16_bit_mixed_signedness_accelerated Bool32
    integer_dot_product_accumulating_saturating32_bit_unsigned_accelerated Bool32
    integer_dot_product_accumulating_saturating32_bit_signed_accelerated Bool32
    integer_dot_product_accumulating_saturating32_bit_mixed_signedness_accelerated Bool32
    integer_dot_product_accumulating_saturating64_bit_unsigned_accelerated Bool32
    integer_dot_product_accumulating_saturating64_bit_signed_accelerated Bool32
    integer_dot_product_accumulating_saturating64_bit_mixed_signedness_accelerated Bool32
} 

// PhysicalDeviceTexelBufferAlignmentProperties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceTexelBufferAlignmentProperties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    storage_texel_buffer_offset_alignment_bytes DeviceSize
    storage_texel_buffer_offset_single_texel_alignment Bool32
    uniform_texel_buffer_offset_alignment_bytes DeviceSize
    uniform_texel_buffer_offset_single_texel_alignment Bool32
} 

// FormatProperties3 extends VkFormatProperties2
pub struct FormatProperties3 {
mut:
    s_type                       StructureType
    p_next                       voidptr
    linear_tiling_features       FormatFeatureFlags2
    optimal_tiling_features      FormatFeatureFlags2
    buffer_features              FormatFeatureFlags2
} 

// PhysicalDeviceMaintenance4Features extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMaintenance4Features {
mut:
    s_type                 StructureType
    p_next                 voidptr
    maintenance4           Bool32
} 

// PhysicalDeviceMaintenance4Properties extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceMaintenance4Properties {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_buffer_size        DeviceSize
} 

pub struct DeviceBufferMemoryRequirements {
mut:
    s_type                           StructureType
    p_next                           voidptr
    p_create_info                    &BufferCreateInfo
} 

pub struct DeviceImageMemoryRequirements {
mut:
    s_type                          StructureType
    p_next                          voidptr
    p_create_info                   &ImageCreateInfo
    plane_aspect                    ImageAspectFlagBits
} 

type VkGetPhysicalDeviceToolProperties = fn (     C.PhysicalDevice,     &u32,     &PhysicalDeviceToolProperties) Result

pub fn get_physical_device_tool_properties(
    physical_device                                 C.PhysicalDevice,
    p_tool_count                                    &u32,
    p_tool_properties                               &PhysicalDeviceToolProperties) Result {
      f := VkGetPhysicalDeviceToolProperties((*loader_p).get_sym('vkGetPhysicalDeviceToolProperties'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceToolProperties': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_tool_count,
    p_tool_properties)
}


type VkCreatePrivateDataSlot = fn (     C.Device,     &PrivateDataSlotCreateInfo,     &AllocationCallbacks,     &C.PrivateDataSlot) Result

pub fn create_private_data_slot(
    device                                          C.Device,
    p_create_info                                   &PrivateDataSlotCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_private_data_slot                             &C.PrivateDataSlot) Result {
      f := VkCreatePrivateDataSlot((*loader_p).get_sym('vkCreatePrivateDataSlot'
    ) or { 
        println("Couldn't load symbol for 'vkCreatePrivateDataSlot': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_private_data_slot)
}


type VkDestroyPrivateDataSlot = fn (     C.Device,     C.PrivateDataSlot,     &AllocationCallbacks) 

pub fn destroy_private_data_slot(
    device                                          C.Device,
    private_data_slot                               C.PrivateDataSlot,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyPrivateDataSlot((*loader_p).get_sym('vkDestroyPrivateDataSlot'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyPrivateDataSlot': ${err}")
        return 
    })
    f(
    device,
    private_data_slot,
    p_allocator)
}


type VkSetPrivateData = fn (     C.Device,     ObjectType,     u64,     C.PrivateDataSlot,     u64) Result

pub fn set_private_data(
    device                                          C.Device,
    object_type                                     ObjectType,
    object_handle                                   u64,
    private_data_slot                               C.PrivateDataSlot,
    data                                            u64) Result {
      f := VkSetPrivateData((*loader_p).get_sym('vkSetPrivateData'
    ) or { 
        println("Couldn't load symbol for 'vkSetPrivateData': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    object_type,
    object_handle,
    private_data_slot,
    data)
}


type VkGetPrivateData = fn (     C.Device,     ObjectType,     u64,     C.PrivateDataSlot,     &u64) 

pub fn get_private_data(
    device                                          C.Device,
    object_type                                     ObjectType,
    object_handle                                   u64,
    private_data_slot                               C.PrivateDataSlot,
    p_data                                          &u64)  {
      f := VkGetPrivateData((*loader_p).get_sym('vkGetPrivateData'
    ) or { 
        println("Couldn't load symbol for 'vkGetPrivateData': ${err}")
        return 
    })
    f(
    device,
    object_type,
    object_handle,
    private_data_slot,
    p_data)
}


type VkCmdSetEvent2 = fn (     C.CommandBuffer,     C.Event,     &DependencyInfo) 

pub fn cmd_set_event2(
    command_buffer                                  C.CommandBuffer,
    event                                           C.Event,
    p_dependency_info                               &DependencyInfo)  {
      f := VkCmdSetEvent2((*loader_p).get_sym('vkCmdSetEvent2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetEvent2': ${err}")
        return 
    })
    f(
    command_buffer,
    event,
    p_dependency_info)
}


type VkCmdResetEvent2 = fn (     C.CommandBuffer,     C.Event,     PipelineStageFlags2) 

pub fn cmd_reset_event2(
    command_buffer                                  C.CommandBuffer,
    event                                           C.Event,
    stage_mask                                      PipelineStageFlags2)  {
      f := VkCmdResetEvent2((*loader_p).get_sym('vkCmdResetEvent2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdResetEvent2': ${err}")
        return 
    })
    f(
    command_buffer,
    event,
    stage_mask)
}


type VkCmdWaitEvents2 = fn (     C.CommandBuffer,     u32,     &C.Event,     &DependencyInfo) 

pub fn cmd_wait_events2(
    command_buffer                                  C.CommandBuffer,
    event_count                                     u32,
    p_events                                        &C.Event,
    p_dependency_infos                              &DependencyInfo)  {
      f := VkCmdWaitEvents2((*loader_p).get_sym('vkCmdWaitEvents2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdWaitEvents2': ${err}")
        return 
    })
    f(
    command_buffer,
    event_count,
    p_events,
    p_dependency_infos)
}


type VkCmdPipelineBarrier2 = fn (     C.CommandBuffer,     &DependencyInfo) 

pub fn cmd_pipeline_barrier2(
    command_buffer                                  C.CommandBuffer,
    p_dependency_info                               &DependencyInfo)  {
      f := VkCmdPipelineBarrier2((*loader_p).get_sym('vkCmdPipelineBarrier2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdPipelineBarrier2': ${err}")
        return 
    })
    f(
    command_buffer,
    p_dependency_info)
}


type VkCmdWriteTimestamp2 = fn (     C.CommandBuffer,     PipelineStageFlags2,     C.QueryPool,     u32) 

pub fn cmd_write_timestamp2(
    command_buffer                                  C.CommandBuffer,
    stage                                           PipelineStageFlags2,
    query_pool                                      C.QueryPool,
    query                                           u32)  {
      f := VkCmdWriteTimestamp2((*loader_p).get_sym('vkCmdWriteTimestamp2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdWriteTimestamp2': ${err}")
        return 
    })
    f(
    command_buffer,
    stage,
    query_pool,
    query)
}


type VkQueueSubmit2 = fn (     C.Queue,     u32,     &SubmitInfo2,     C.Fence) Result

pub fn queue_submit2(
    queue                                           C.Queue,
    submit_count                                    u32,
    p_submits                                       &SubmitInfo2,
    fence                                           C.Fence) Result {
      f := VkQueueSubmit2((*loader_p).get_sym('vkQueueSubmit2'
    ) or { 
        println("Couldn't load symbol for 'vkQueueSubmit2': ${err}")
        return Result.error_unknown
    })
    return f(
    queue,
    submit_count,
    p_submits,
    fence)
}


type VkCmdCopyBuffer2 = fn (     C.CommandBuffer,     &CopyBufferInfo2) 

pub fn cmd_copy_buffer2(
    command_buffer                                  C.CommandBuffer,
    p_copy_buffer_info                              &CopyBufferInfo2)  {
      f := VkCmdCopyBuffer2((*loader_p).get_sym('vkCmdCopyBuffer2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyBuffer2': ${err}")
        return 
    })
    f(
    command_buffer,
    p_copy_buffer_info)
}


type VkCmdCopyImage2 = fn (     C.CommandBuffer,     &CopyImageInfo2) 

pub fn cmd_copy_image2(
    command_buffer                                  C.CommandBuffer,
    p_copy_image_info                               &CopyImageInfo2)  {
      f := VkCmdCopyImage2((*loader_p).get_sym('vkCmdCopyImage2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyImage2': ${err}")
        return 
    })
    f(
    command_buffer,
    p_copy_image_info)
}


type VkCmdCopyBufferToImage2 = fn (     C.CommandBuffer,     &CopyBufferToImageInfo2) 

pub fn cmd_copy_buffer_to_image2(
    command_buffer                                  C.CommandBuffer,
    p_copy_buffer_to_image_info                     &CopyBufferToImageInfo2)  {
      f := VkCmdCopyBufferToImage2((*loader_p).get_sym('vkCmdCopyBufferToImage2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyBufferToImage2': ${err}")
        return 
    })
    f(
    command_buffer,
    p_copy_buffer_to_image_info)
}


type VkCmdCopyImageToBuffer2 = fn (     C.CommandBuffer,     &CopyImageToBufferInfo2) 

pub fn cmd_copy_image_to_buffer2(
    command_buffer                                  C.CommandBuffer,
    p_copy_image_to_buffer_info                     &CopyImageToBufferInfo2)  {
      f := VkCmdCopyImageToBuffer2((*loader_p).get_sym('vkCmdCopyImageToBuffer2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyImageToBuffer2': ${err}")
        return 
    })
    f(
    command_buffer,
    p_copy_image_to_buffer_info)
}


type VkCmdBlitImage2 = fn (     C.CommandBuffer,     &BlitImageInfo2) 

pub fn cmd_blit_image2(
    command_buffer                                  C.CommandBuffer,
    p_blit_image_info                               &BlitImageInfo2)  {
      f := VkCmdBlitImage2((*loader_p).get_sym('vkCmdBlitImage2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBlitImage2': ${err}")
        return 
    })
    f(
    command_buffer,
    p_blit_image_info)
}


type VkCmdResolveImage2 = fn (     C.CommandBuffer,     &ResolveImageInfo2) 

pub fn cmd_resolve_image2(
    command_buffer                                  C.CommandBuffer,
    p_resolve_image_info                            &ResolveImageInfo2)  {
      f := VkCmdResolveImage2((*loader_p).get_sym('vkCmdResolveImage2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdResolveImage2': ${err}")
        return 
    })
    f(
    command_buffer,
    p_resolve_image_info)
}


type VkCmdBeginRendering = fn (     C.CommandBuffer,     &RenderingInfo) 

pub fn cmd_begin_rendering(
    command_buffer                                  C.CommandBuffer,
    p_rendering_info                                &RenderingInfo)  {
      f := VkCmdBeginRendering((*loader_p).get_sym('vkCmdBeginRendering'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBeginRendering': ${err}")
        return 
    })
    f(
    command_buffer,
    p_rendering_info)
}


type VkCmdEndRendering = fn (     C.CommandBuffer) 

pub fn cmd_end_rendering(
    command_buffer                                  C.CommandBuffer)  {
      f := VkCmdEndRendering((*loader_p).get_sym('vkCmdEndRendering'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEndRendering': ${err}")
        return 
    })
    f(
    command_buffer)
}


type VkCmdSetCullMode = fn (     C.CommandBuffer,     CullModeFlags) 

pub fn cmd_set_cull_mode(
    command_buffer                                  C.CommandBuffer,
    cull_mode                                       CullModeFlags)  {
      f := VkCmdSetCullMode((*loader_p).get_sym('vkCmdSetCullMode'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetCullMode': ${err}")
        return 
    })
    f(
    command_buffer,
    cull_mode)
}


type VkCmdSetFrontFace = fn (     C.CommandBuffer,     FrontFace) 

pub fn cmd_set_front_face(
    command_buffer                                  C.CommandBuffer,
    front_face                                      FrontFace)  {
      f := VkCmdSetFrontFace((*loader_p).get_sym('vkCmdSetFrontFace'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetFrontFace': ${err}")
        return 
    })
    f(
    command_buffer,
    front_face)
}


type VkCmdSetPrimitiveTopology = fn (     C.CommandBuffer,     PrimitiveTopology) 

pub fn cmd_set_primitive_topology(
    command_buffer                                  C.CommandBuffer,
    primitive_topology                              PrimitiveTopology)  {
      f := VkCmdSetPrimitiveTopology((*loader_p).get_sym('vkCmdSetPrimitiveTopology'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetPrimitiveTopology': ${err}")
        return 
    })
    f(
    command_buffer,
    primitive_topology)
}


type VkCmdSetViewportWithCount = fn (     C.CommandBuffer,     u32,     &Viewport) 

pub fn cmd_set_viewport_with_count(
    command_buffer                                  C.CommandBuffer,
    viewport_count                                  u32,
    p_viewports                                     &Viewport)  {
      f := VkCmdSetViewportWithCount((*loader_p).get_sym('vkCmdSetViewportWithCount'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetViewportWithCount': ${err}")
        return 
    })
    f(
    command_buffer,
    viewport_count,
    p_viewports)
}


type VkCmdSetScissorWithCount = fn (     C.CommandBuffer,     u32,     &Rect2D) 

pub fn cmd_set_scissor_with_count(
    command_buffer                                  C.CommandBuffer,
    scissor_count                                   u32,
    p_scissors                                      &Rect2D)  {
      f := VkCmdSetScissorWithCount((*loader_p).get_sym('vkCmdSetScissorWithCount'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetScissorWithCount': ${err}")
        return 
    })
    f(
    command_buffer,
    scissor_count,
    p_scissors)
}


type VkCmdBindVertexBuffers2 = fn (     C.CommandBuffer,     u32,     u32,     &C.Buffer,     &DeviceSize,     &DeviceSize,     &DeviceSize) 

pub fn cmd_bind_vertex_buffers2(
    command_buffer                                  C.CommandBuffer,
    first_binding                                   u32,
    binding_count                                   u32,
    p_buffers                                       &C.Buffer,
    p_offsets                                       &DeviceSize,
    p_sizes                                         &DeviceSize,
    p_strides                                       &DeviceSize)  {
      f := VkCmdBindVertexBuffers2((*loader_p).get_sym('vkCmdBindVertexBuffers2'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindVertexBuffers2': ${err}")
        return 
    })
    f(
    command_buffer,
    first_binding,
    binding_count,
    p_buffers,
    p_offsets,
    p_sizes,
    p_strides)
}


type VkCmdSetDepthTestEnable = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_depth_test_enable(
    command_buffer                                  C.CommandBuffer,
    depth_test_enable                               Bool32)  {
      f := VkCmdSetDepthTestEnable((*loader_p).get_sym('vkCmdSetDepthTestEnable'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthTestEnable': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_test_enable)
}


type VkCmdSetDepthWriteEnable = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_depth_write_enable(
    command_buffer                                  C.CommandBuffer,
    depth_write_enable                              Bool32)  {
      f := VkCmdSetDepthWriteEnable((*loader_p).get_sym('vkCmdSetDepthWriteEnable'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthWriteEnable': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_write_enable)
}


type VkCmdSetDepthCompareOp = fn (     C.CommandBuffer,     CompareOp) 

pub fn cmd_set_depth_compare_op(
    command_buffer                                  C.CommandBuffer,
    depth_compare_op                                CompareOp)  {
      f := VkCmdSetDepthCompareOp((*loader_p).get_sym('vkCmdSetDepthCompareOp'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthCompareOp': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_compare_op)
}


type VkCmdSetDepthBoundsTestEnable = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_depth_bounds_test_enable(
    command_buffer                                  C.CommandBuffer,
    depth_bounds_test_enable                        Bool32)  {
      f := VkCmdSetDepthBoundsTestEnable((*loader_p).get_sym('vkCmdSetDepthBoundsTestEnable'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthBoundsTestEnable': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_bounds_test_enable)
}


type VkCmdSetStencilTestEnable = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_stencil_test_enable(
    command_buffer                                  C.CommandBuffer,
    stencil_test_enable                             Bool32)  {
      f := VkCmdSetStencilTestEnable((*loader_p).get_sym('vkCmdSetStencilTestEnable'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetStencilTestEnable': ${err}")
        return 
    })
    f(
    command_buffer,
    stencil_test_enable)
}


type VkCmdSetStencilOp = fn (     C.CommandBuffer,     StencilFaceFlags,     StencilOp,     StencilOp,     StencilOp,     CompareOp) 

pub fn cmd_set_stencil_op(
    command_buffer                                  C.CommandBuffer,
    face_mask                                       StencilFaceFlags,
    fail_op                                         StencilOp,
    pass_op                                         StencilOp,
    depth_fail_op                                   StencilOp,
    compare_op                                      CompareOp)  {
      f := VkCmdSetStencilOp((*loader_p).get_sym('vkCmdSetStencilOp'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetStencilOp': ${err}")
        return 
    })
    f(
    command_buffer,
    face_mask,
    fail_op,
    pass_op,
    depth_fail_op,
    compare_op)
}


type VkCmdSetRasterizerDiscardEnable = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_rasterizer_discard_enable(
    command_buffer                                  C.CommandBuffer,
    rasterizer_discard_enable                       Bool32)  {
      f := VkCmdSetRasterizerDiscardEnable((*loader_p).get_sym('vkCmdSetRasterizerDiscardEnable'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetRasterizerDiscardEnable': ${err}")
        return 
    })
    f(
    command_buffer,
    rasterizer_discard_enable)
}


type VkCmdSetDepthBiasEnable = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_depth_bias_enable(
    command_buffer                                  C.CommandBuffer,
    depth_bias_enable                               Bool32)  {
      f := VkCmdSetDepthBiasEnable((*loader_p).get_sym('vkCmdSetDepthBiasEnable'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthBiasEnable': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_bias_enable)
}


type VkCmdSetPrimitiveRestartEnable = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_primitive_restart_enable(
    command_buffer                                  C.CommandBuffer,
    primitive_restart_enable                        Bool32)  {
      f := VkCmdSetPrimitiveRestartEnable((*loader_p).get_sym('vkCmdSetPrimitiveRestartEnable'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetPrimitiveRestartEnable': ${err}")
        return 
    })
    f(
    command_buffer,
    primitive_restart_enable)
}


type VkGetDeviceBufferMemoryRequirements = fn (     C.Device,     &DeviceBufferMemoryRequirements,     &MemoryRequirements2) 

pub fn get_device_buffer_memory_requirements(
    device                                          C.Device,
    p_info                                          &DeviceBufferMemoryRequirements,
    p_memory_requirements                           &MemoryRequirements2)  {
      f := VkGetDeviceBufferMemoryRequirements((*loader_p).get_sym('vkGetDeviceBufferMemoryRequirements'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceBufferMemoryRequirements': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_memory_requirements)
}


type VkGetDeviceImageMemoryRequirements = fn (     C.Device,     &DeviceImageMemoryRequirements,     &MemoryRequirements2) 

pub fn get_device_image_memory_requirements(
    device                                          C.Device,
    p_info                                          &DeviceImageMemoryRequirements,
    p_memory_requirements                           &MemoryRequirements2)  {
      f := VkGetDeviceImageMemoryRequirements((*loader_p).get_sym('vkGetDeviceImageMemoryRequirements'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceImageMemoryRequirements': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_memory_requirements)
}


type VkGetDeviceImageSparseMemoryRequirements = fn (     C.Device,     &DeviceImageMemoryRequirements,     &u32,     &SparseImageMemoryRequirements2) 

pub fn get_device_image_sparse_memory_requirements(
    device                                          C.Device,
    p_info                                          &DeviceImageMemoryRequirements,
    p_sparse_memory_requirement_count               &u32,
    p_sparse_memory_requirements                    &SparseImageMemoryRequirements2)  {
      f := VkGetDeviceImageSparseMemoryRequirements((*loader_p).get_sym('vkGetDeviceImageSparseMemoryRequirements'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceImageSparseMemoryRequirements': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_sparse_memory_requirement_count,
    p_sparse_memory_requirements)
}




// VK_KHR_surface is a preprocessor guard. Do not pass it to API calls.
const khr_surface = 1
pub type C.SurfaceKHR = voidptr
pub const khr_surface_spec_version          = 25
pub const khr_surface_extension_name        = "VK_KHR_surface"

pub enum PresentModeKHR {
    present_mode_immediate_khr = int(0)
    present_mode_mailbox_khr = int(1)
    present_mode_fifo_khr = int(2)
    present_mode_fifo_relaxed_khr = int(3)
    present_mode_shared_demand_refresh_khr = int(1000111000)
    present_mode_shared_continuous_refresh_khr = int(1000111001)
    present_mode_max_enum_khr = int(0x7FFFFFFF)
}


pub enum ColorSpaceKHR {
    color_space_srgb_nonlinear_khr = int(0)
    color_space_display_p3_nonlinear_ext = int(1000104001)
    color_space_extended_srgb_linear_ext = int(1000104002)
    color_space_display_p3_linear_ext = int(1000104003)
    color_space_dci_p3_nonlinear_ext = int(1000104004)
    color_space_bt709_linear_ext = int(1000104005)
    color_space_bt709_nonlinear_ext = int(1000104006)
    color_space_bt2020_linear_ext = int(1000104007)
    color_space_hdr10_st2084_ext = int(1000104008)
    color_space_dolbyvision_ext = int(1000104009)
    color_space_hdr10_hlg_ext = int(1000104010)
    color_space_adobergb_linear_ext = int(1000104011)
    color_space_adobergb_nonlinear_ext = int(1000104012)
    color_space_pass_through_ext = int(1000104013)
    color_space_extended_srgb_nonlinear_ext = int(1000104014)
    color_space_display_native_amd = int(1000213000)
    color_space_max_enum_khr = int(0x7FFFFFFF)
}


pub enum SurfaceTransformFlagBitsKHR {
    surface_transform_identity_bit_khr = int(0x00000001)
    surface_transform_rotate_90_bit_khr = int(0x00000002)
    surface_transform_rotate_180_bit_khr = int(0x00000004)
    surface_transform_rotate_270_bit_khr = int(0x00000008)
    surface_transform_horizontal_mirror_bit_khr = int(0x00000010)
    surface_transform_horizontal_mirror_rotate_90_bit_khr = int(0x00000020)
    surface_transform_horizontal_mirror_rotate_180_bit_khr = int(0x00000040)
    surface_transform_horizontal_mirror_rotate_270_bit_khr = int(0x00000080)
    surface_transform_inherit_bit_khr = int(0x00000100)
    surface_transform_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}


pub enum CompositeAlphaFlagBitsKHR {
    composite_alpha_opaque_bit_khr = int(0x00000001)
    composite_alpha_pre_multiplied_bit_khr = int(0x00000002)
    composite_alpha_post_multiplied_bit_khr = int(0x00000004)
    composite_alpha_inherit_bit_khr = int(0x00000008)
    composite_alpha_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type CompositeAlphaFlagsKHR = u32
pub type SurfaceTransformFlagsKHR = u32
pub struct SurfaceCapabilitiesKHR {
mut:
    min_image_count                      u32
    max_image_count                      u32
    current_extent                       Extent2D
    min_image_extent                     Extent2D
    max_image_extent                     Extent2D
    max_image_array_layers               u32
    supported_transforms                 SurfaceTransformFlagsKHR
    current_transform                    SurfaceTransformFlagBitsKHR
    supported_composite_alpha            CompositeAlphaFlagsKHR
    supported_usage_flags                ImageUsageFlags
} 

pub struct SurfaceFormatKHR {
mut:
    format                 Format
    color_space            ColorSpaceKHR
} 

type VkDestroySurfaceKHR = fn (     C.Instance,     C.SurfaceKHR,     &AllocationCallbacks) 

pub fn destroy_surface_khr(
    instance                                        C.Instance,
    surface                                         C.SurfaceKHR,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroySurfaceKHR((*loader_p).get_sym('vkDestroySurfaceKHR'
    ) or { 
        println("Couldn't load symbol for 'vkDestroySurfaceKHR': ${err}")
        return 
    })
    f(
    instance,
    surface,
    p_allocator)
}


type VkGetPhysicalDeviceSurfaceSupportKHR = fn (     C.PhysicalDevice,     u32,     C.SurfaceKHR,     &Bool32) Result

pub fn get_physical_device_surface_support_khr(
    physical_device                                 C.PhysicalDevice,
    queue_family_index                              u32,
    surface                                         C.SurfaceKHR,
    p_supported                                     &Bool32) Result {
      f := VkGetPhysicalDeviceSurfaceSupportKHR((*loader_p).get_sym('vkGetPhysicalDeviceSurfaceSupportKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSurfaceSupportKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    queue_family_index,
    surface,
    p_supported)
}


type VkGetPhysicalDeviceSurfaceCapabilitiesKHR = fn (     C.PhysicalDevice,     C.SurfaceKHR,     &SurfaceCapabilitiesKHR) Result

pub fn get_physical_device_surface_capabilities_khr(
    physical_device                                 C.PhysicalDevice,
    surface                                         C.SurfaceKHR,
    p_surface_capabilities                          &SurfaceCapabilitiesKHR) Result {
      f := VkGetPhysicalDeviceSurfaceCapabilitiesKHR((*loader_p).get_sym('vkGetPhysicalDeviceSurfaceCapabilitiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSurfaceCapabilitiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    surface,
    p_surface_capabilities)
}


type VkGetPhysicalDeviceSurfaceFormatsKHR = fn (     C.PhysicalDevice,     C.SurfaceKHR,     &u32,     &SurfaceFormatKHR) Result

pub fn get_physical_device_surface_formats_khr(
    physical_device                                 C.PhysicalDevice,
    surface                                         C.SurfaceKHR,
    p_surface_format_count                          &u32,
    p_surface_formats                               &SurfaceFormatKHR) Result {
      f := VkGetPhysicalDeviceSurfaceFormatsKHR((*loader_p).get_sym('vkGetPhysicalDeviceSurfaceFormatsKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSurfaceFormatsKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    surface,
    p_surface_format_count,
    p_surface_formats)
}


type VkGetPhysicalDeviceSurfacePresentModesKHR = fn (     C.PhysicalDevice,     C.SurfaceKHR,     &u32,     &PresentModeKHR) Result

pub fn get_physical_device_surface_present_modes_khr(
    physical_device                                 C.PhysicalDevice,
    surface                                         C.SurfaceKHR,
    p_present_mode_count                            &u32,
    p_present_modes                                 &PresentModeKHR) Result {
      f := VkGetPhysicalDeviceSurfacePresentModesKHR((*loader_p).get_sym('vkGetPhysicalDeviceSurfacePresentModesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSurfacePresentModesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    surface,
    p_present_mode_count,
    p_present_modes)
}




// VK_KHR_swapchain is a preprocessor guard. Do not pass it to API calls.
const khr_swapchain = 1
pub type C.SwapchainKHR = voidptr
pub const khr_swapchain_spec_version        = 70
pub const khr_swapchain_extension_name      = "VK_KHR_swapchain"

pub enum SwapchainCreateFlagBitsKHR {
    swapchain_create_split_instance_bind_regions_bit_khr = int(0x00000001)
    swapchain_create_protected_bit_khr = int(0x00000002)
    swapchain_create_mutable_format_bit_khr = int(0x00000004)
    swapchain_create_deferred_memory_allocation_bit_ext = int(0x00000008)
    swapchain_create_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type SwapchainCreateFlagsKHR = u32

pub enum DeviceGroupPresentModeFlagBitsKHR {
    device_group_present_mode_local_bit_khr = int(0x00000001)
    device_group_present_mode_remote_bit_khr = int(0x00000002)
    device_group_present_mode_sum_bit_khr = int(0x00000004)
    device_group_present_mode_local_multi_device_bit_khr = int(0x00000008)
    device_group_present_mode_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type DeviceGroupPresentModeFlagsKHR = u32
pub struct SwapchainCreateInfoKHR {
mut:
    s_type                               StructureType
    p_next                               voidptr
    flags                                SwapchainCreateFlagsKHR
    surface                              C.SurfaceKHR
    min_image_count                      u32
    image_format                         Format
    image_color_space                    ColorSpaceKHR
    image_extent                         Extent2D
    image_array_layers                   u32
    image_usage                          ImageUsageFlags
    image_sharing_mode                   SharingMode
    queue_family_index_count             u32
    p_queue_family_indices               &u32
    pre_transform                        SurfaceTransformFlagBitsKHR
    composite_alpha                      CompositeAlphaFlagBitsKHR
    present_mode                         PresentModeKHR
    clipped                              Bool32
    old_swapchain                        C.SwapchainKHR
} 

pub struct PresentInfoKHR {
mut:
    s_type                       StructureType
    p_next                       voidptr
    wait_semaphore_count         u32
    p_wait_semaphores            &C.Semaphore
    swapchain_count              u32
    p_swapchains                 &C.SwapchainKHR
    p_image_indices              &u32
    p_results                    &Result
} 

// ImageSwapchainCreateInfoKHR extends VkImageCreateInfo
pub struct ImageSwapchainCreateInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    swapchain              C.SwapchainKHR
} 

// BindImageMemorySwapchainInfoKHR extends VkBindImageMemoryInfo
pub struct BindImageMemorySwapchainInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    swapchain              C.SwapchainKHR
    image_index            u32
} 

pub struct AcquireNextImageInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    swapchain              C.SwapchainKHR
    timeout                u64
    semaphore              C.Semaphore
    fence                  C.Fence
    device_mask            u32
} 

pub struct DeviceGroupPresentCapabilitiesKHR {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    present_mask                            []u32
    modes                                   DeviceGroupPresentModeFlagsKHR
} 

// DeviceGroupPresentInfoKHR extends VkPresentInfoKHR
pub struct DeviceGroupPresentInfoKHR {
mut:
    s_type                                     StructureType
    p_next                                     voidptr
    swapchain_count                            u32
    p_device_masks                             &u32
    mode                                       DeviceGroupPresentModeFlagBitsKHR
} 

// DeviceGroupSwapchainCreateInfoKHR extends VkSwapchainCreateInfoKHR
pub struct DeviceGroupSwapchainCreateInfoKHR {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    modes                                   DeviceGroupPresentModeFlagsKHR
} 

type VkCreateSwapchainKHR = fn (     C.Device,     &SwapchainCreateInfoKHR,     &AllocationCallbacks,     &C.SwapchainKHR) Result

pub fn create_swapchain_khr(
    device                                          C.Device,
    p_create_info                                   &SwapchainCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_swapchain                                     &C.SwapchainKHR) Result {
      f := VkCreateSwapchainKHR((*loader_p).get_sym('vkCreateSwapchainKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateSwapchainKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_swapchain)
}


type VkDestroySwapchainKHR = fn (     C.Device,     C.SwapchainKHR,     &AllocationCallbacks) 

pub fn destroy_swapchain_khr(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroySwapchainKHR((*loader_p).get_sym('vkDestroySwapchainKHR'
    ) or { 
        println("Couldn't load symbol for 'vkDestroySwapchainKHR': ${err}")
        return 
    })
    f(
    device,
    swapchain,
    p_allocator)
}


type VkGetSwapchainImagesKHR = fn (     C.Device,     C.SwapchainKHR,     &u32,     &C.Image) Result

pub fn get_swapchain_images_khr(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR,
    p_swapchain_image_count                         &u32,
    p_swapchain_images                              &C.Image) Result {
      f := VkGetSwapchainImagesKHR((*loader_p).get_sym('vkGetSwapchainImagesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetSwapchainImagesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain,
    p_swapchain_image_count,
    p_swapchain_images)
}


type VkAcquireNextImageKHR = fn (     C.Device,     C.SwapchainKHR,     u64,     C.Semaphore,     C.Fence,     &u32) Result

pub fn acquire_next_image_khr(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR,
    timeout                                         u64,
    semaphore                                       C.Semaphore,
    fence                                           C.Fence,
    p_image_index                                   &u32) Result {
      f := VkAcquireNextImageKHR((*loader_p).get_sym('vkAcquireNextImageKHR'
    ) or { 
        println("Couldn't load symbol for 'vkAcquireNextImageKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain,
    timeout,
    semaphore,
    fence,
    p_image_index)
}


type VkQueuePresentKHR = fn (     C.Queue,     &PresentInfoKHR) Result

pub fn queue_present_khr(
    queue                                           C.Queue,
    p_present_info                                  &PresentInfoKHR) Result {
      f := VkQueuePresentKHR((*loader_p).get_sym('vkQueuePresentKHR'
    ) or { 
        println("Couldn't load symbol for 'vkQueuePresentKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    queue,
    p_present_info)
}


type VkGetDeviceGroupPresentCapabilitiesKHR = fn (     C.Device,     &DeviceGroupPresentCapabilitiesKHR) Result

pub fn get_device_group_present_capabilities_khr(
    device                                          C.Device,
    p_device_group_present_capabilities             &DeviceGroupPresentCapabilitiesKHR) Result {
      f := VkGetDeviceGroupPresentCapabilitiesKHR((*loader_p).get_sym('vkGetDeviceGroupPresentCapabilitiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceGroupPresentCapabilitiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_device_group_present_capabilities)
}


type VkGetDeviceGroupSurfacePresentModesKHR = fn (     C.Device,     C.SurfaceKHR,     &DeviceGroupPresentModeFlagsKHR) Result

pub fn get_device_group_surface_present_modes_khr(
    device                                          C.Device,
    surface                                         C.SurfaceKHR,
    p_modes                                         &DeviceGroupPresentModeFlagsKHR) Result {
      f := VkGetDeviceGroupSurfacePresentModesKHR((*loader_p).get_sym('vkGetDeviceGroupSurfacePresentModesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceGroupSurfacePresentModesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    surface,
    p_modes)
}


type VkGetPhysicalDevicePresentRectanglesKHR = fn (     C.PhysicalDevice,     C.SurfaceKHR,     &u32,     &Rect2D) Result

pub fn get_physical_device_present_rectangles_khr(
    physical_device                                 C.PhysicalDevice,
    surface                                         C.SurfaceKHR,
    p_rect_count                                    &u32,
    p_rects                                         &Rect2D) Result {
      f := VkGetPhysicalDevicePresentRectanglesKHR((*loader_p).get_sym('vkGetPhysicalDevicePresentRectanglesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDevicePresentRectanglesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    surface,
    p_rect_count,
    p_rects)
}


type VkAcquireNextImage2KHR = fn (     C.Device,     &AcquireNextImageInfoKHR,     &u32) Result

pub fn acquire_next_image2_khr(
    device                                          C.Device,
    p_acquire_info                                  &AcquireNextImageInfoKHR,
    p_image_index                                   &u32) Result {
      f := VkAcquireNextImage2KHR((*loader_p).get_sym('vkAcquireNextImage2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkAcquireNextImage2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_acquire_info,
    p_image_index)
}




// VK_KHR_display is a preprocessor guard. Do not pass it to API calls.
const khr_display = 1
pub type C.DisplayKHR = voidptr
pub type C.DisplayModeKHR = voidptr
pub const khr_display_spec_version          = 23
pub const khr_display_extension_name        = "VK_KHR_display"
pub type DisplayModeCreateFlagsKHR = u32

pub enum DisplayPlaneAlphaFlagBitsKHR {
    display_plane_alpha_opaque_bit_khr = int(0x00000001)
    display_plane_alpha_global_bit_khr = int(0x00000002)
    display_plane_alpha_per_pixel_bit_khr = int(0x00000004)
    display_plane_alpha_per_pixel_premultiplied_bit_khr = int(0x00000008)
    display_plane_alpha_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type DisplayPlaneAlphaFlagsKHR = u32
pub type DisplaySurfaceCreateFlagsKHR = u32
pub struct DisplayModeParametersKHR {
mut:
    visible_region    Extent2D
    refresh_rate      u32
} 

pub struct DisplayModeCreateInfoKHR {
mut:
    s_type                             StructureType
    p_next                             voidptr
    flags                              DisplayModeCreateFlagsKHR
    parameters                         DisplayModeParametersKHR
} 

pub struct DisplayModePropertiesKHR {
mut:
    display_mode                      C.DisplayModeKHR
    parameters                        DisplayModeParametersKHR
} 

pub struct DisplayPlaneCapabilitiesKHR {
mut:
    supported_alpha                    DisplayPlaneAlphaFlagsKHR
    min_src_position                   Offset2D
    max_src_position                   Offset2D
    min_src_extent                     Extent2D
    max_src_extent                     Extent2D
    min_dst_position                   Offset2D
    max_dst_position                   Offset2D
    min_dst_extent                     Extent2D
    max_dst_extent                     Extent2D
} 

pub struct DisplayPlanePropertiesKHR {
mut:
    current_display     C.DisplayKHR
    current_stack_index u32
} 

pub struct DisplayPropertiesKHR {
mut:
    display                           C.DisplayKHR
    display_name                      &char
    physical_dimensions               Extent2D
    physical_resolution               Extent2D
    supported_transforms              SurfaceTransformFlagsKHR
    plane_reorder_possible            Bool32
    persistent_content                Bool32
} 

pub struct DisplaySurfaceCreateInfoKHR {
mut:
    s_type                                StructureType
    p_next                                voidptr
    flags                                 DisplaySurfaceCreateFlagsKHR
    display_mode                          C.DisplayModeKHR
    plane_index                           u32
    plane_stack_index                     u32
    transform                             SurfaceTransformFlagBitsKHR
    global_alpha                          f32
    alpha_mode                            DisplayPlaneAlphaFlagBitsKHR
    image_extent                          Extent2D
} 

type VkGetPhysicalDeviceDisplayPropertiesKHR = fn (     C.PhysicalDevice,     &u32,     &DisplayPropertiesKHR) Result

pub fn get_physical_device_display_properties_khr(
    physical_device                                 C.PhysicalDevice,
    p_property_count                                &u32,
    p_properties                                    &DisplayPropertiesKHR) Result {
      f := VkGetPhysicalDeviceDisplayPropertiesKHR((*loader_p).get_sym('vkGetPhysicalDeviceDisplayPropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceDisplayPropertiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_property_count,
    p_properties)
}


type VkGetPhysicalDeviceDisplayPlanePropertiesKHR = fn (     C.PhysicalDevice,     &u32,     &DisplayPlanePropertiesKHR) Result

pub fn get_physical_device_display_plane_properties_khr(
    physical_device                                 C.PhysicalDevice,
    p_property_count                                &u32,
    p_properties                                    &DisplayPlanePropertiesKHR) Result {
      f := VkGetPhysicalDeviceDisplayPlanePropertiesKHR((*loader_p).get_sym('vkGetPhysicalDeviceDisplayPlanePropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceDisplayPlanePropertiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_property_count,
    p_properties)
}


type VkGetDisplayPlaneSupportedDisplaysKHR = fn (     C.PhysicalDevice,     u32,     &u32,     &C.DisplayKHR) Result

pub fn get_display_plane_supported_displays_khr(
    physical_device                                 C.PhysicalDevice,
    plane_index                                     u32,
    p_display_count                                 &u32,
    p_displays                                      &C.DisplayKHR) Result {
      f := VkGetDisplayPlaneSupportedDisplaysKHR((*loader_p).get_sym('vkGetDisplayPlaneSupportedDisplaysKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDisplayPlaneSupportedDisplaysKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    plane_index,
    p_display_count,
    p_displays)
}


type VkGetDisplayModePropertiesKHR = fn (     C.PhysicalDevice,     C.DisplayKHR,     &u32,     &DisplayModePropertiesKHR) Result

pub fn get_display_mode_properties_khr(
    physical_device                                 C.PhysicalDevice,
    display                                         C.DisplayKHR,
    p_property_count                                &u32,
    p_properties                                    &DisplayModePropertiesKHR) Result {
      f := VkGetDisplayModePropertiesKHR((*loader_p).get_sym('vkGetDisplayModePropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDisplayModePropertiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    display,
    p_property_count,
    p_properties)
}


type VkCreateDisplayModeKHR = fn (     C.PhysicalDevice,     C.DisplayKHR,     &DisplayModeCreateInfoKHR,     &AllocationCallbacks,     &C.DisplayModeKHR) Result

pub fn create_display_mode_khr(
    physical_device                                 C.PhysicalDevice,
    display                                         C.DisplayKHR,
    p_create_info                                   &DisplayModeCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_mode                                          &C.DisplayModeKHR) Result {
      f := VkCreateDisplayModeKHR((*loader_p).get_sym('vkCreateDisplayModeKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateDisplayModeKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    display,
    p_create_info,
    p_allocator,
    p_mode)
}


type VkGetDisplayPlaneCapabilitiesKHR = fn (     C.PhysicalDevice,     C.DisplayModeKHR,     u32,     &DisplayPlaneCapabilitiesKHR) Result

pub fn get_display_plane_capabilities_khr(
    physical_device                                 C.PhysicalDevice,
    mode                                            C.DisplayModeKHR,
    plane_index                                     u32,
    p_capabilities                                  &DisplayPlaneCapabilitiesKHR) Result {
      f := VkGetDisplayPlaneCapabilitiesKHR((*loader_p).get_sym('vkGetDisplayPlaneCapabilitiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDisplayPlaneCapabilitiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    mode,
    plane_index,
    p_capabilities)
}


type VkCreateDisplayPlaneSurfaceKHR = fn (     C.Instance,     &DisplaySurfaceCreateInfoKHR,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_display_plane_surface_khr(
    instance                                        C.Instance,
    p_create_info                                   &DisplaySurfaceCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateDisplayPlaneSurfaceKHR((*loader_p).get_sym('vkCreateDisplayPlaneSurfaceKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateDisplayPlaneSurfaceKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}




// VK_KHR_display_swapchain is a preprocessor guard. Do not pass it to API calls.
const khr_display_swapchain = 1
pub const khr_display_swapchain_spec_version = 10
pub const khr_display_swapchain_extension_name = "VK_KHR_display_swapchain"
// DisplayPresentInfoKHR extends VkPresentInfoKHR
pub struct DisplayPresentInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    src_rect               Rect2D
    dst_rect               Rect2D
    persistent             Bool32
} 

type VkCreateSharedSwapchainsKHR = fn (     C.Device,     u32,     &SwapchainCreateInfoKHR,     &AllocationCallbacks,     &C.SwapchainKHR) Result

pub fn create_shared_swapchains_khr(
    device                                          C.Device,
    swapchain_count                                 u32,
    p_create_infos                                  &SwapchainCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_swapchains                                    &C.SwapchainKHR) Result {
      f := VkCreateSharedSwapchainsKHR((*loader_p).get_sym('vkCreateSharedSwapchainsKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateSharedSwapchainsKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain_count,
    p_create_infos,
    p_allocator,
    p_swapchains)
}




// VK_KHR_xlib_surface is a preprocessor guard. Do not pass it to API calls.
const khr_xlib_surface = 1
pub const khr_xlib_surface_spec_version     = 6
pub const khr_xlib_surface_extension_name   = "VK_KHR_xlib_surface"
pub type XlibSurfaceCreateFlagsKHR = u32
pub struct XlibSurfaceCreateInfoKHR {
mut:
    s_type                             StructureType
    p_next                             voidptr
    flags                              XlibSurfaceCreateFlagsKHR
    dpy                                &C.DisplayKHR
    window                             voidptr
} 

type VkCreateXlibSurfaceKHR = fn (     C.Instance,     &XlibSurfaceCreateInfoKHR,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_xlib_surface_khr(
    instance                                        C.Instance,
    p_create_info                                   &XlibSurfaceCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateXlibSurfaceKHR((*loader_p).get_sym('vkCreateXlibSurfaceKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateXlibSurfaceKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}


type VkGetPhysicalDeviceXlibPresentationSupportKHR = fn (     C.PhysicalDevice,     u32,     &C.DisplayKHR,     voidptr) Bool32

pub fn get_physical_device_xlib_presentation_support_khr(
    physical_device                                 C.PhysicalDevice,
    queue_family_index                              u32,
    dpy                                             &C.DisplayKHR,
    visual_id                                       voidptr) Bool32 {
      f := VkGetPhysicalDeviceXlibPresentationSupportKHR((*loader_p).get_sym("vkGetPhysicalDeviceXlibPresentationSupportKHR"
    ) or { 
        panic("Couldn't load symbol for 'vkGetPhysicalDeviceXlibPresentationSupportKHR': ${err}") })
    return f(
    physical_device,
    queue_family_index,
    dpy,
    visual_id)
}




// VK_KHR_xcb_surface is a preprocessor guard. Do not pass it to API calls.
const khr_xcb_surface = 1
pub const khr_xcb_surface_spec_version      = 6
pub const khr_xcb_surface_extension_name    = "VK_KHR_xcb_surface"
pub type XcbSurfaceCreateFlagsKHR = u32
pub struct XcbSurfaceCreateInfoKHR {
mut:
    s_type                            StructureType
    p_next                            voidptr
    flags                             XcbSurfaceCreateFlagsKHR
    connection                        voidptr
    window                            voidptr
} 

type VkCreateXcbSurfaceKHR = fn (     C.Instance,     &XcbSurfaceCreateInfoKHR,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_xcb_surface_khr(
    instance                                        C.Instance,
    p_create_info                                   &XcbSurfaceCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateXcbSurfaceKHR((*loader_p).get_sym('vkCreateXcbSurfaceKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateXcbSurfaceKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}


type VkGetPhysicalDeviceXcbPresentationSupportKHR = fn (     C.PhysicalDevice,     u32,     voidptr,     voidptr) Bool32

pub fn get_physical_device_xcb_presentation_support_khr(
    physical_device                                 C.PhysicalDevice,
    queue_family_index                              u32,
    connection                                      voidptr,
    visual_id                                       voidptr) Bool32 {
      f := VkGetPhysicalDeviceXcbPresentationSupportKHR((*loader_p).get_sym("vkGetPhysicalDeviceXcbPresentationSupportKHR"
    ) or { 
        panic("Couldn't load symbol for 'vkGetPhysicalDeviceXcbPresentationSupportKHR': ${err}") })
    return f(
    physical_device,
    queue_family_index,
    connection,
    visual_id)
}




// VK_KHR_wayland_surface is a preprocessor guard. Do not pass it to API calls.
const khr_wayland_surface = 1
pub const khr_wayland_surface_spec_version  = 6
pub const khr_wayland_surface_extension_name = "VK_KHR_wayland_surface"
pub type WaylandSurfaceCreateFlagsKHR = u32
pub struct WaylandSurfaceCreateInfoKHR {
mut:
    s_type                                StructureType
    p_next                                voidptr
    flags                                 WaylandSurfaceCreateFlagsKHR
    display                               voidptr
    surface                               voidptr
} 

type VkCreateWaylandSurfaceKHR = fn (     C.Instance,     &WaylandSurfaceCreateInfoKHR,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_wayland_surface_khr(
    instance                                        C.Instance,
    p_create_info                                   &WaylandSurfaceCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateWaylandSurfaceKHR((*loader_p).get_sym('vkCreateWaylandSurfaceKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateWaylandSurfaceKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}


type VkGetPhysicalDeviceWaylandPresentationSupportKHR = fn (     C.PhysicalDevice,     u32,     voidptr) Bool32

pub fn get_physical_device_wayland_presentation_support_khr(
    physical_device                                 C.PhysicalDevice,
    queue_family_index                              u32,
    display                                         voidptr) Bool32 {
      f := VkGetPhysicalDeviceWaylandPresentationSupportKHR((*loader_p).get_sym("vkGetPhysicalDeviceWaylandPresentationSupportKHR"
    ) or { 
        panic("Couldn't load symbol for 'vkGetPhysicalDeviceWaylandPresentationSupportKHR': ${err}") })
    return f(
    physical_device,
    queue_family_index,
    display)
}




// VK_KHR_android_surface is a preprocessor guard. Do not pass it to API calls.
const khr_android_surface = 1
pub const khr_android_surface_spec_version  = 6
pub const khr_android_surface_extension_name = "VK_KHR_android_surface"
pub type AndroidSurfaceCreateFlagsKHR = u32
pub struct AndroidSurfaceCreateInfoKHR {
mut:
    s_type                                StructureType
    p_next                                voidptr
    flags                                 AndroidSurfaceCreateFlagsKHR
    window                                voidptr
} 

type VkCreateAndroidSurfaceKHR = fn (     C.Instance,     &AndroidSurfaceCreateInfoKHR,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_android_surface_khr(
    instance                                        C.Instance,
    p_create_info                                   &AndroidSurfaceCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateAndroidSurfaceKHR((*loader_p).get_sym('vkCreateAndroidSurfaceKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateAndroidSurfaceKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}




// VK_KHR_win32_surface is a preprocessor guard. Do not pass it to API calls.
const khr_win32_surface = 1
pub const khr_win32_surface_spec_version    = 6
pub const khr_win32_surface_extension_name  = "VK_KHR_win32_surface"
pub type Win32SurfaceCreateFlagsKHR = u32
pub struct Win32SurfaceCreateInfoKHR {
mut:
    s_type                              StructureType
    p_next                              voidptr
    flags                               Win32SurfaceCreateFlagsKHR
    hinstance                           voidptr
    hwnd                                voidptr
} 

type VkCreateWin32SurfaceKHR = fn (     C.Instance,     &Win32SurfaceCreateInfoKHR,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_win32_surface_khr(
    instance                                        C.Instance,
    p_create_info                                   &Win32SurfaceCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateWin32SurfaceKHR((*loader_p).get_sym('vkCreateWin32SurfaceKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateWin32SurfaceKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}


type VkGetPhysicalDeviceWin32PresentationSupportKHR = fn (     C.PhysicalDevice,     u32) Bool32

pub fn get_physical_device_win32_presentation_support_khr(
    physical_device                                 C.PhysicalDevice,
    queue_family_index                              u32) Bool32 {
      f := VkGetPhysicalDeviceWin32PresentationSupportKHR((*loader_p).get_sym("vkGetPhysicalDeviceWin32PresentationSupportKHR"
    ) or { 
        panic("Couldn't load symbol for 'vkGetPhysicalDeviceWin32PresentationSupportKHR': ${err}") })
    return f(
    physical_device,
    queue_family_index)
}




// VK_KHR_sampler_mirror_clamp_to_edge is a preprocessor guard. Do not pass it to API calls.
const khr_sampler_mirror_clamp_to_edge = 1
pub const khr_sampler_mirror_clamp_to_edge_spec_version = 3
pub const khr_sampler_mirror_clamp_to_edge_extension_name = "VK_KHR_sampler_mirror_clamp_to_edge"


// VK_KHR_video_queue is a preprocessor guard. Do not pass it to API calls.
const khr_video_queue = 1
pub type C.VideoSessionKHR = voidptr
pub type C.VideoSessionParametersKHR = voidptr
pub const khr_video_queue_spec_version      = 8
pub const khr_video_queue_extension_name    = "VK_KHR_video_queue"

pub enum QueryResultStatusKHR {
    query_result_status_error_khr = int(-1)
    query_result_status_not_ready_khr = int(0)
    query_result_status_complete_khr = int(1)
    query_result_status_insufficient_bitstream_buffer_range_khr = int(-1000299000)
    query_result_status_max_enum_khr = int(0x7FFFFFFF)
}


pub enum VideoCodecOperationFlagBitsKHR {
    video_codec_operation_none_khr = int(0)
    video_codec_operation_decode_h264_bit_khr = int(0x00000001)
    video_codec_operation_decode_h265_bit_khr = int(0x00000002)
    video_codec_operation_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoCodecOperationFlagsKHR = u32

pub enum VideoChromaSubsamplingFlagBitsKHR {
    video_chroma_subsampling_invalid_khr = int(0)
    video_chroma_subsampling_monochrome_bit_khr = int(0x00000001)
    video_chroma_subsampling_420_bit_khr = int(0x00000002)
    video_chroma_subsampling_422_bit_khr = int(0x00000004)
    video_chroma_subsampling_444_bit_khr = int(0x00000008)
    video_chroma_subsampling_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoChromaSubsamplingFlagsKHR = u32

pub enum VideoComponentBitDepthFlagBitsKHR {
    video_component_bit_depth_invalid_khr = int(0)
    video_component_bit_depth_8_bit_khr = int(0x00000001)
    video_component_bit_depth_10_bit_khr = int(0x00000004)
    video_component_bit_depth_12_bit_khr = int(0x00000010)
    video_component_bit_depth_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoComponentBitDepthFlagsKHR = u32

pub enum VideoCapabilityFlagBitsKHR {
    video_capability_protected_content_bit_khr = int(0x00000001)
    video_capability_separate_reference_images_bit_khr = int(0x00000002)
    video_capability_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoCapabilityFlagsKHR = u32

pub enum VideoSessionCreateFlagBitsKHR {
    video_session_create_protected_content_bit_khr = int(0x00000001)
    video_session_create_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoSessionCreateFlagsKHR = u32
pub type VideoSessionParametersCreateFlagsKHR = u32
pub type VideoBeginCodingFlagsKHR = u32
pub type VideoEndCodingFlagsKHR = u32

pub enum VideoCodingControlFlagBitsKHR {
    video_coding_control_reset_bit_khr = int(0x00000001)
    video_coding_control_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoCodingControlFlagsKHR = u32
// QueueFamilyQueryResultStatusPropertiesKHR extends VkQueueFamilyProperties2
pub struct QueueFamilyQueryResultStatusPropertiesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    query_result_status_support Bool32
} 

// QueueFamilyVideoPropertiesKHR extends VkQueueFamilyProperties2
pub struct QueueFamilyVideoPropertiesKHR {
mut:
    s_type                               StructureType
    p_next                               voidptr
    video_codec_operations               VideoCodecOperationFlagsKHR
} 

// VideoProfileInfoKHR extends VkQueryPoolCreateInfo
pub struct VideoProfileInfoKHR {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    video_codec_operation                   VideoCodecOperationFlagBitsKHR
    chroma_subsampling                      VideoChromaSubsamplingFlagsKHR
    luma_bit_depth                          VideoComponentBitDepthFlagsKHR
    chroma_bit_depth                        VideoComponentBitDepthFlagsKHR
} 

// VideoProfileListInfoKHR extends VkPhysicalDeviceImageFormatInfo2,VkPhysicalDeviceVideoFormatInfoKHR,VkImageCreateInfo,VkBufferCreateInfo
pub struct VideoProfileListInfoKHR {
mut:
    s_type                              StructureType
    p_next                              voidptr
    profile_count                       u32
    p_profiles                          &VideoProfileInfoKHR
} 

pub struct VideoCapabilitiesKHR {
mut:
    s_type                           StructureType
    p_next                           voidptr
    flags                            VideoCapabilityFlagsKHR
    min_bitstream_buffer_offset_alignment DeviceSize
    min_bitstream_buffer_size_alignment DeviceSize
    picture_access_granularity       Extent2D
    min_coded_extent                 Extent2D
    max_coded_extent                 Extent2D
    max_dpb_slots                    u32
    max_active_reference_pictures    u32
    std_header_version               ExtensionProperties
} 

pub struct PhysicalDeviceVideoFormatInfoKHR {
mut:
    s_type                   StructureType
    p_next                   voidptr
    image_usage              ImageUsageFlags
} 

pub struct VideoFormatPropertiesKHR {
mut:
    s_type                    StructureType
    p_next                    voidptr
    format                    Format
    component_mapping         ComponentMapping
    image_create_flags        ImageCreateFlags
    image_type                ImageType
    image_tiling              ImageTiling
    image_usage_flags         ImageUsageFlags
} 

pub struct VideoPictureResourceInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    coded_offset           Offset2D
    coded_extent           Extent2D
    base_array_layer       u32
    image_view_binding     C.ImageView
} 

pub struct VideoReferenceSlotInfoKHR {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    slot_index                                  i32
    p_picture_resource                          &VideoPictureResourceInfoKHR
} 

pub struct VideoSessionMemoryRequirementsKHR {
mut:
    s_type                      StructureType
    p_next                      voidptr
    memory_bind_index           u32
    memory_requirements         MemoryRequirements
} 

pub struct BindVideoSessionMemoryInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    memory_bind_index      u32
    memory                 C.DeviceMemory
    memory_offset          DeviceSize
    memory_size            DeviceSize
} 

pub struct VideoSessionCreateInfoKHR {
mut:
    s_type                              StructureType
    p_next                              voidptr
    queue_family_index                  u32
    flags                               VideoSessionCreateFlagsKHR
    p_video_profile                     &VideoProfileInfoKHR
    picture_format                      Format
    max_coded_extent                    Extent2D
    reference_picture_format            Format
    max_dpb_slots                       u32
    max_active_reference_pictures       u32
    p_std_header_version                &ExtensionProperties
} 

pub struct VideoSessionParametersCreateInfoKHR {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    flags                                         VideoSessionParametersCreateFlagsKHR
    video_session_parameters_template             C.VideoSessionParametersKHR
    video_session                                 C.VideoSessionKHR
} 

pub struct VideoSessionParametersUpdateInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    update_sequence_count  u32
} 

pub struct VideoBeginCodingInfoKHR {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    flags                                     VideoBeginCodingFlagsKHR
    video_session                             C.VideoSessionKHR
    video_session_parameters                  C.VideoSessionParametersKHR
    reference_slot_count                      u32
    p_reference_slots                         &VideoReferenceSlotInfoKHR
} 

pub struct VideoEndCodingInfoKHR {
mut:
    s_type                          StructureType
    p_next                          voidptr
    flags                           VideoEndCodingFlagsKHR
} 

pub struct VideoCodingControlInfoKHR {
mut:
    s_type                              StructureType
    p_next                              voidptr
    flags                               VideoCodingControlFlagsKHR
} 

type VkGetPhysicalDeviceVideoCapabilitiesKHR = fn (     C.PhysicalDevice,     &VideoProfileInfoKHR,     &VideoCapabilitiesKHR) Result

pub fn get_physical_device_video_capabilities_khr(
    physical_device                                 C.PhysicalDevice,
    p_video_profile                                 &VideoProfileInfoKHR,
    p_capabilities                                  &VideoCapabilitiesKHR) Result {
      f := VkGetPhysicalDeviceVideoCapabilitiesKHR((*loader_p).get_sym('vkGetPhysicalDeviceVideoCapabilitiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceVideoCapabilitiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_video_profile,
    p_capabilities)
}


type VkGetPhysicalDeviceVideoFormatPropertiesKHR = fn (     C.PhysicalDevice,     &PhysicalDeviceVideoFormatInfoKHR,     &u32,     &VideoFormatPropertiesKHR) Result

pub fn get_physical_device_video_format_properties_khr(
    physical_device                                 C.PhysicalDevice,
    p_video_format_info                             &PhysicalDeviceVideoFormatInfoKHR,
    p_video_format_property_count                   &u32,
    p_video_format_properties                       &VideoFormatPropertiesKHR) Result {
      f := VkGetPhysicalDeviceVideoFormatPropertiesKHR((*loader_p).get_sym('vkGetPhysicalDeviceVideoFormatPropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceVideoFormatPropertiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_video_format_info,
    p_video_format_property_count,
    p_video_format_properties)
}


type VkCreateVideoSessionKHR = fn (     C.Device,     &VideoSessionCreateInfoKHR,     &AllocationCallbacks,     &C.VideoSessionKHR) Result

pub fn create_video_session_khr(
    device                                          C.Device,
    p_create_info                                   &VideoSessionCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_video_session                                 &C.VideoSessionKHR) Result {
      f := VkCreateVideoSessionKHR((*loader_p).get_sym('vkCreateVideoSessionKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateVideoSessionKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_video_session)
}


type VkDestroyVideoSessionKHR = fn (     C.Device,     C.VideoSessionKHR,     &AllocationCallbacks) 

pub fn destroy_video_session_khr(
    device                                          C.Device,
    video_session                                   C.VideoSessionKHR,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyVideoSessionKHR((*loader_p).get_sym('vkDestroyVideoSessionKHR'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyVideoSessionKHR': ${err}")
        return 
    })
    f(
    device,
    video_session,
    p_allocator)
}


type VkGetVideoSessionMemoryRequirementsKHR = fn (     C.Device,     C.VideoSessionKHR,     &u32,     &VideoSessionMemoryRequirementsKHR) Result

pub fn get_video_session_memory_requirements_khr(
    device                                          C.Device,
    video_session                                   C.VideoSessionKHR,
    p_memory_requirements_count                     &u32,
    p_memory_requirements                           &VideoSessionMemoryRequirementsKHR) Result {
      f := VkGetVideoSessionMemoryRequirementsKHR((*loader_p).get_sym('vkGetVideoSessionMemoryRequirementsKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetVideoSessionMemoryRequirementsKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    video_session,
    p_memory_requirements_count,
    p_memory_requirements)
}


type VkBindVideoSessionMemoryKHR = fn (     C.Device,     C.VideoSessionKHR,     u32,     &BindVideoSessionMemoryInfoKHR) Result

pub fn bind_video_session_memory_khr(
    device                                          C.Device,
    video_session                                   C.VideoSessionKHR,
    bind_session_memory_info_count                  u32,
    p_bind_session_memory_infos                     &BindVideoSessionMemoryInfoKHR) Result {
      f := VkBindVideoSessionMemoryKHR((*loader_p).get_sym('vkBindVideoSessionMemoryKHR'
    ) or { 
        println("Couldn't load symbol for 'vkBindVideoSessionMemoryKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    video_session,
    bind_session_memory_info_count,
    p_bind_session_memory_infos)
}


type VkCreateVideoSessionParametersKHR = fn (     C.Device,     &VideoSessionParametersCreateInfoKHR,     &AllocationCallbacks,     &C.VideoSessionParametersKHR) Result

pub fn create_video_session_parameters_khr(
    device                                          C.Device,
    p_create_info                                   &VideoSessionParametersCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_video_session_parameters                      &C.VideoSessionParametersKHR) Result {
      f := VkCreateVideoSessionParametersKHR((*loader_p).get_sym('vkCreateVideoSessionParametersKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateVideoSessionParametersKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_video_session_parameters)
}


type VkUpdateVideoSessionParametersKHR = fn (     C.Device,     C.VideoSessionParametersKHR,     &VideoSessionParametersUpdateInfoKHR) Result

pub fn update_video_session_parameters_khr(
    device                                          C.Device,
    video_session_parameters                        C.VideoSessionParametersKHR,
    p_update_info                                   &VideoSessionParametersUpdateInfoKHR) Result {
      f := VkUpdateVideoSessionParametersKHR((*loader_p).get_sym('vkUpdateVideoSessionParametersKHR'
    ) or { 
        println("Couldn't load symbol for 'vkUpdateVideoSessionParametersKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    video_session_parameters,
    p_update_info)
}


type VkDestroyVideoSessionParametersKHR = fn (     C.Device,     C.VideoSessionParametersKHR,     &AllocationCallbacks) 

pub fn destroy_video_session_parameters_khr(
    device                                          C.Device,
    video_session_parameters                        C.VideoSessionParametersKHR,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyVideoSessionParametersKHR((*loader_p).get_sym('vkDestroyVideoSessionParametersKHR'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyVideoSessionParametersKHR': ${err}")
        return 
    })
    f(
    device,
    video_session_parameters,
    p_allocator)
}


type VkCmdBeginVideoCodingKHR = fn (     C.CommandBuffer,     &VideoBeginCodingInfoKHR) 

pub fn cmd_begin_video_coding_khr(
    command_buffer                                  C.CommandBuffer,
    p_begin_info                                    &VideoBeginCodingInfoKHR)  {
      f := VkCmdBeginVideoCodingKHR((*loader_p).get_sym('vkCmdBeginVideoCodingKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBeginVideoCodingKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_begin_info)
}


type VkCmdEndVideoCodingKHR = fn (     C.CommandBuffer,     &VideoEndCodingInfoKHR) 

pub fn cmd_end_video_coding_khr(
    command_buffer                                  C.CommandBuffer,
    p_end_coding_info                               &VideoEndCodingInfoKHR)  {
      f := VkCmdEndVideoCodingKHR((*loader_p).get_sym('vkCmdEndVideoCodingKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEndVideoCodingKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_end_coding_info)
}


type VkCmdControlVideoCodingKHR = fn (     C.CommandBuffer,     &VideoCodingControlInfoKHR) 

pub fn cmd_control_video_coding_khr(
    command_buffer                                  C.CommandBuffer,
    p_coding_control_info                           &VideoCodingControlInfoKHR)  {
      f := VkCmdControlVideoCodingKHR((*loader_p).get_sym('vkCmdControlVideoCodingKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdControlVideoCodingKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_coding_control_info)
}




// VK_KHR_video_decode_queue is a preprocessor guard. Do not pass it to API calls.
const khr_video_decode_queue = 1
pub const khr_video_decode_queue_spec_version = 7
pub const khr_video_decode_queue_extension_name = "VK_KHR_video_decode_queue"

pub enum VideoDecodeCapabilityFlagBitsKHR {
    video_decode_capability_dpb_and_output_coincide_bit_khr = int(0x00000001)
    video_decode_capability_dpb_and_output_distinct_bit_khr = int(0x00000002)
    video_decode_capability_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoDecodeCapabilityFlagsKHR = u32

pub enum VideoDecodeUsageFlagBitsKHR {
    video_decode_usage_default_khr = int(0)
    video_decode_usage_transcoding_bit_khr = int(0x00000001)
    video_decode_usage_offline_bit_khr = int(0x00000002)
    video_decode_usage_streaming_bit_khr = int(0x00000004)
    video_decode_usage_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoDecodeUsageFlagsKHR = u32
pub type VideoDecodeFlagsKHR = u32
// VideoDecodeCapabilitiesKHR extends VkVideoCapabilitiesKHR
pub struct VideoDecodeCapabilitiesKHR {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    flags                                  VideoDecodeCapabilityFlagsKHR
} 

// VideoDecodeUsageInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub struct VideoDecodeUsageInfoKHR {
mut:
    s_type                            StructureType
    p_next                            voidptr
    video_usage_hints                 VideoDecodeUsageFlagsKHR
} 

pub struct VideoDecodeInfoKHR {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    flags                                     VideoDecodeFlagsKHR
    src_buffer                                C.Buffer
    src_buffer_offset                         DeviceSize
    src_buffer_range                          DeviceSize
    dst_picture_resource                      VideoPictureResourceInfoKHR
    p_setup_reference_slot                    &VideoReferenceSlotInfoKHR
    reference_slot_count                      u32
    p_reference_slots                         &VideoReferenceSlotInfoKHR
} 

type VkCmdDecodeVideoKHR = fn (     C.CommandBuffer,     &VideoDecodeInfoKHR) 

pub fn cmd_decode_video_khr(
    command_buffer                                  C.CommandBuffer,
    p_decode_info                                   &VideoDecodeInfoKHR)  {
      f := VkCmdDecodeVideoKHR((*loader_p).get_sym('vkCmdDecodeVideoKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDecodeVideoKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_decode_info)
}




// VK_KHR_video_decode_h264 is a preprocessor guard. Do not pass it to API calls.
const khr_video_decode_h264 = 1
pub const khr_video_decode_h264_spec_version = 8
pub const khr_video_decode_h264_extension_name = "VK_KHR_video_decode_h264"

pub enum VideoDecodeH264PictureLayoutFlagBitsKHR {
    video_decode_h264_picture_layout_progressive_khr = int(0)
    video_decode_h264_picture_layout_interlaced_interleaved_lines_bit_khr = int(0x00000001)
    video_decode_h264_picture_layout_interlaced_separate_planes_bit_khr = int(0x00000002)
    video_decode_h264_picture_layout_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoDecodeH264PictureLayoutFlagsKHR = u32
// VideoDecodeH264ProfileInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub struct VideoDecodeH264ProfileInfoKHR {
mut:
    s_type                                           StructureType
    p_next                                           voidptr
    std_profile_idc                                  C.StdVideoH264ProfileIdc
    picture_layout                                   VideoDecodeH264PictureLayoutFlagBitsKHR
} 

// VideoDecodeH264CapabilitiesKHR extends VkVideoCapabilitiesKHR
pub struct VideoDecodeH264CapabilitiesKHR {
mut:
    s_type                      StructureType
    p_next                      voidptr
    max_level_idc               C.StdVideoH264LevelIdc
    field_offset_granularity    Offset2D
} 

// VideoDecodeH264SessionParametersAddInfoKHR extends VkVideoSessionParametersUpdateInfoKHR
pub struct VideoDecodeH264SessionParametersAddInfoKHR {
mut:
    s_type                                         StructureType
    p_next                                         voidptr
    std_sps_count                                  u32
    p_std_sp_ss                                    &C.StdVideoH264SequenceParameterSet
    std_pps_count                                  u32
    p_std_pp_ss                                    &C.StdVideoH264PictureParameterSet
} 

// VideoDecodeH264SessionParametersCreateInfoKHR extends VkVideoSessionParametersCreateInfoKHR
pub struct VideoDecodeH264SessionParametersCreateInfoKHR {
mut:
    s_type                                                     StructureType
    p_next                                                     voidptr
    max_std_sps_count                                          u32
    max_std_pps_count                                          u32
    p_parameters_add_info                                      &VideoDecodeH264SessionParametersAddInfoKHR
} 

// VideoDecodeH264PictureInfoKHR extends VkVideoDecodeInfoKHR
pub struct VideoDecodeH264PictureInfoKHR {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    p_std_picture_info                          &C.StdVideoDecodeH264PictureInfo
    slice_count                                 u32
    p_slice_offsets                             &u32
} 

// VideoDecodeH264DpbSlotInfoKHR extends VkVideoReferenceSlotInfoKHR
pub struct VideoDecodeH264DpbSlotInfoKHR {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    p_std_reference_info                          &C.StdVideoDecodeH264ReferenceInfo
} 



// VK_KHR_dynamic_rendering is a preprocessor guard. Do not pass it to API calls.
const khr_dynamic_rendering = 1
pub const khr_dynamic_rendering_spec_version = 1
pub const khr_dynamic_rendering_extension_name = "VK_KHR_dynamic_rendering"
pub type RenderingFlagBitsKHR = RenderingFlagBits

pub type RenderingInfoKHR = RenderingInfo

pub type RenderingAttachmentInfoKHR = RenderingAttachmentInfo

pub type PipelineRenderingCreateInfoKHR = PipelineRenderingCreateInfo

pub type PhysicalDeviceDynamicRenderingFeaturesKHR = PhysicalDeviceDynamicRenderingFeatures

pub type CommandBufferInheritanceRenderingInfoKHR = CommandBufferInheritanceRenderingInfo

// RenderingFragmentShadingRateAttachmentInfoKHR extends VkRenderingInfo
pub struct RenderingFragmentShadingRateAttachmentInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image_view             C.ImageView
    image_layout           ImageLayout
    shading_rate_attachment_texel_size Extent2D
} 

// RenderingFragmentDensityMapAttachmentInfoEXT extends VkRenderingInfo
pub struct RenderingFragmentDensityMapAttachmentInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image_view             C.ImageView
    image_layout           ImageLayout
} 

// AttachmentSampleCountInfoAMD extends VkCommandBufferInheritanceInfo,VkGraphicsPipelineCreateInfo
pub struct AttachmentSampleCountInfoAMD {
mut:
    s_type                              StructureType
    p_next                              voidptr
    color_attachment_count              u32
    p_color_attachment_samples          &SampleCountFlagBits
    depth_stencil_attachment_samples    SampleCountFlagBits
} 

pub type AttachmentSampleCountInfoNV = AttachmentSampleCountInfoAMD

// MultiviewPerViewAttributesInfoNVX extends VkCommandBufferInheritanceInfo,VkGraphicsPipelineCreateInfo,VkRenderingInfo
pub struct MultiviewPerViewAttributesInfoNVX {
mut:
    s_type                 StructureType
    p_next                 voidptr
    per_view_attributes    Bool32
    per_view_attributes_position_x_only Bool32
} 

type VkCmdBeginRenderingKHR = fn (     C.CommandBuffer,     &RenderingInfo) 

pub fn cmd_begin_rendering_khr(
    command_buffer                                  C.CommandBuffer,
    p_rendering_info                                &RenderingInfo)  {
      f := VkCmdBeginRenderingKHR((*loader_p).get_sym('vkCmdBeginRenderingKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBeginRenderingKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_rendering_info)
}


type VkCmdEndRenderingKHR = fn (     C.CommandBuffer) 

pub fn cmd_end_rendering_khr(
    command_buffer                                  C.CommandBuffer)  {
      f := VkCmdEndRenderingKHR((*loader_p).get_sym('vkCmdEndRenderingKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEndRenderingKHR': ${err}")
        return 
    })
    f(
    command_buffer)
}




// VK_KHR_multiview is a preprocessor guard. Do not pass it to API calls.
const khr_multiview = 1
pub const khr_multiview_spec_version        = 1
pub const khr_multiview_extension_name      = "VK_KHR_multiview"
pub type RenderPassMultiviewCreateInfoKHR = RenderPassMultiviewCreateInfo

pub type PhysicalDeviceMultiviewFeaturesKHR = PhysicalDeviceMultiviewFeatures

pub type PhysicalDeviceMultiviewPropertiesKHR = PhysicalDeviceMultiviewProperties



// VK_KHR_get_physical_device_properties2 is a preprocessor guard. Do not pass it to API calls.
const khr_get_physical_device_properties2 = 1
pub const khr_get_physical_device_properties_2_spec_version = 2
pub const khr_get_physical_device_properties_2_extension_name = "VK_KHR_get_physical_device_properties2"
pub type PhysicalDeviceFeatures2KHR = PhysicalDeviceFeatures2

pub type PhysicalDeviceProperties2KHR = PhysicalDeviceProperties2

pub type FormatProperties2KHR = FormatProperties2

pub type ImageFormatProperties2KHR = ImageFormatProperties2

pub type PhysicalDeviceImageFormatInfo2KHR = PhysicalDeviceImageFormatInfo2

pub type QueueFamilyProperties2KHR = QueueFamilyProperties2

pub type PhysicalDeviceMemoryProperties2KHR = PhysicalDeviceMemoryProperties2

pub type SparseImageFormatProperties2KHR = SparseImageFormatProperties2

pub type PhysicalDeviceSparseImageFormatInfo2KHR = PhysicalDeviceSparseImageFormatInfo2

type VkGetPhysicalDeviceFeatures2KHR = fn (     C.PhysicalDevice,     &PhysicalDeviceFeatures2) 

pub fn get_physical_device_features2_khr(
    physical_device                                 C.PhysicalDevice,
    p_features                                      &PhysicalDeviceFeatures2)  {
      f := VkGetPhysicalDeviceFeatures2KHR((*loader_p).get_sym('vkGetPhysicalDeviceFeatures2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceFeatures2KHR': ${err}")
        return 
    })
    f(
    physical_device,
    p_features)
}


type VkGetPhysicalDeviceProperties2KHR = fn (     C.PhysicalDevice,     &PhysicalDeviceProperties2) 

pub fn get_physical_device_properties2_khr(
    physical_device                                 C.PhysicalDevice,
    p_properties                                    &PhysicalDeviceProperties2)  {
      f := VkGetPhysicalDeviceProperties2KHR((*loader_p).get_sym('vkGetPhysicalDeviceProperties2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceProperties2KHR': ${err}")
        return 
    })
    f(
    physical_device,
    p_properties)
}


type VkGetPhysicalDeviceFormatProperties2KHR = fn (     C.PhysicalDevice,     Format,     &FormatProperties2) 

pub fn get_physical_device_format_properties2_khr(
    physical_device                                 C.PhysicalDevice,
    format                                          Format,
    p_format_properties                             &FormatProperties2)  {
      f := VkGetPhysicalDeviceFormatProperties2KHR((*loader_p).get_sym('vkGetPhysicalDeviceFormatProperties2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceFormatProperties2KHR': ${err}")
        return 
    })
    f(
    physical_device,
    format,
    p_format_properties)
}


type VkGetPhysicalDeviceImageFormatProperties2KHR = fn (     C.PhysicalDevice,     &PhysicalDeviceImageFormatInfo2,     &ImageFormatProperties2) Result

pub fn get_physical_device_image_format_properties2_khr(
    physical_device                                 C.PhysicalDevice,
    p_image_format_info                             &PhysicalDeviceImageFormatInfo2,
    p_image_format_properties                       &ImageFormatProperties2) Result {
      f := VkGetPhysicalDeviceImageFormatProperties2KHR((*loader_p).get_sym('vkGetPhysicalDeviceImageFormatProperties2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceImageFormatProperties2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_image_format_info,
    p_image_format_properties)
}


type VkGetPhysicalDeviceQueueFamilyProperties2KHR = fn (     C.PhysicalDevice,     &u32,     &QueueFamilyProperties2) 

pub fn get_physical_device_queue_family_properties2_khr(
    physical_device                                 C.PhysicalDevice,
    p_queue_family_property_count                   &u32,
    p_queue_family_properties                       &QueueFamilyProperties2)  {
      f := VkGetPhysicalDeviceQueueFamilyProperties2KHR((*loader_p).get_sym('vkGetPhysicalDeviceQueueFamilyProperties2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceQueueFamilyProperties2KHR': ${err}")
        return 
    })
    f(
    physical_device,
    p_queue_family_property_count,
    p_queue_family_properties)
}


type VkGetPhysicalDeviceMemoryProperties2KHR = fn (     C.PhysicalDevice,     &PhysicalDeviceMemoryProperties2) 

pub fn get_physical_device_memory_properties2_khr(
    physical_device                                 C.PhysicalDevice,
    p_memory_properties                             &PhysicalDeviceMemoryProperties2)  {
      f := VkGetPhysicalDeviceMemoryProperties2KHR((*loader_p).get_sym('vkGetPhysicalDeviceMemoryProperties2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceMemoryProperties2KHR': ${err}")
        return 
    })
    f(
    physical_device,
    p_memory_properties)
}


type VkGetPhysicalDeviceSparseImageFormatProperties2KHR = fn (     C.PhysicalDevice,     &PhysicalDeviceSparseImageFormatInfo2,     &u32,     &SparseImageFormatProperties2) 

pub fn get_physical_device_sparse_image_format_properties2_khr(
    physical_device                                 C.PhysicalDevice,
    p_format_info                                   &PhysicalDeviceSparseImageFormatInfo2,
    p_property_count                                &u32,
    p_properties                                    &SparseImageFormatProperties2)  {
      f := VkGetPhysicalDeviceSparseImageFormatProperties2KHR((*loader_p).get_sym('vkGetPhysicalDeviceSparseImageFormatProperties2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSparseImageFormatProperties2KHR': ${err}")
        return 
    })
    f(
    physical_device,
    p_format_info,
    p_property_count,
    p_properties)
}




// VK_KHR_device_group is a preprocessor guard. Do not pass it to API calls.
const khr_device_group = 1
pub const khr_device_group_spec_version     = 4
pub const khr_device_group_extension_name   = "VK_KHR_device_group"
pub type PeerMemoryFeatureFlagBitsKHR = PeerMemoryFeatureFlagBits

pub type MemoryAllocateFlagBitsKHR = MemoryAllocateFlagBits

pub type MemoryAllocateFlagsInfoKHR = MemoryAllocateFlagsInfo

pub type DeviceGroupRenderPassBeginInfoKHR = DeviceGroupRenderPassBeginInfo

pub type DeviceGroupCommandBufferBeginInfoKHR = DeviceGroupCommandBufferBeginInfo

pub type DeviceGroupSubmitInfoKHR = DeviceGroupSubmitInfo

pub type DeviceGroupBindSparseInfoKHR = DeviceGroupBindSparseInfo

pub type BindBufferMemoryDeviceGroupInfoKHR = BindBufferMemoryDeviceGroupInfo

pub type BindImageMemoryDeviceGroupInfoKHR = BindImageMemoryDeviceGroupInfo

type VkGetDeviceGroupPeerMemoryFeaturesKHR = fn (     C.Device,     u32,     u32,     u32,     &PeerMemoryFeatureFlags) 

pub fn get_device_group_peer_memory_features_khr(
    device                                          C.Device,
    heap_index                                      u32,
    local_device_index                              u32,
    remote_device_index                             u32,
    p_peer_memory_features                          &PeerMemoryFeatureFlags)  {
      f := VkGetDeviceGroupPeerMemoryFeaturesKHR((*loader_p).get_sym('vkGetDeviceGroupPeerMemoryFeaturesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceGroupPeerMemoryFeaturesKHR': ${err}")
        return 
    })
    f(
    device,
    heap_index,
    local_device_index,
    remote_device_index,
    p_peer_memory_features)
}


type VkCmdSetDeviceMaskKHR = fn (     C.CommandBuffer,     u32) 

pub fn cmd_set_device_mask_khr(
    command_buffer                                  C.CommandBuffer,
    device_mask                                     u32)  {
      f := VkCmdSetDeviceMaskKHR((*loader_p).get_sym('vkCmdSetDeviceMaskKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDeviceMaskKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    device_mask)
}


type VkCmdDispatchBaseKHR = fn (     C.CommandBuffer,     u32,     u32,     u32,     u32,     u32,     u32) 

pub fn cmd_dispatch_base_khr(
    command_buffer                                  C.CommandBuffer,
    base_group_x                                    u32,
    base_group_y                                    u32,
    base_group_z                                    u32,
    group_count_x                                   u32,
    group_count_y                                   u32,
    group_count_z                                   u32)  {
      f := VkCmdDispatchBaseKHR((*loader_p).get_sym('vkCmdDispatchBaseKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDispatchBaseKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    base_group_x,
    base_group_y,
    base_group_z,
    group_count_x,
    group_count_y,
    group_count_z)
}




// VK_KHR_shader_draw_parameters is a preprocessor guard. Do not pass it to API calls.
const khr_shader_draw_parameters = 1
pub const khr_shader_draw_parameters_spec_version = 1
pub const khr_shader_draw_parameters_extension_name = "VK_KHR_shader_draw_parameters"


// VK_KHR_maintenance1 is a preprocessor guard. Do not pass it to API calls.
const khr_maintenance1 = 1
pub const khr_maintenance_1_spec_version    = 2
pub const khr_maintenance_1_extension_name  = "VK_KHR_maintenance1"
pub const khr_maintenance1_spec_version     = khr_maintenance_1_spec_version
pub const khr_maintenance1_extension_name   = khr_maintenance_1_extension_name
type VkTrimCommandPoolKHR = fn (     C.Device,     C.CommandPool,     CommandPoolTrimFlags) 

pub fn trim_command_pool_khr(
    device                                          C.Device,
    command_pool                                    C.CommandPool,
    flags                                           CommandPoolTrimFlags)  {
      f := VkTrimCommandPoolKHR((*loader_p).get_sym('vkTrimCommandPoolKHR'
    ) or { 
        println("Couldn't load symbol for 'vkTrimCommandPoolKHR': ${err}")
        return 
    })
    f(
    device,
    command_pool,
    flags)
}




// VK_KHR_device_group_creation is a preprocessor guard. Do not pass it to API calls.
const khr_device_group_creation = 1
pub const khr_device_group_creation_spec_version = 1
pub const khr_device_group_creation_extension_name = "VK_KHR_device_group_creation"
pub const max_device_group_size_khr         = max_device_group_size
pub type PhysicalDeviceGroupPropertiesKHR = PhysicalDeviceGroupProperties

pub type DeviceGroupDeviceCreateInfoKHR = DeviceGroupDeviceCreateInfo

type VkEnumeratePhysicalDeviceGroupsKHR = fn (     C.Instance,     &u32,     &PhysicalDeviceGroupProperties) Result

pub fn enumerate_physical_device_groups_khr(
    instance                                        C.Instance,
    p_physical_device_group_count                   &u32,
    p_physical_device_group_properties              &PhysicalDeviceGroupProperties) Result {
      f := VkEnumeratePhysicalDeviceGroupsKHR((*loader_p).get_sym('vkEnumeratePhysicalDeviceGroupsKHR'
    ) or { 
        println("Couldn't load symbol for 'vkEnumeratePhysicalDeviceGroupsKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_physical_device_group_count,
    p_physical_device_group_properties)
}




// VK_KHR_external_memory_capabilities is a preprocessor guard. Do not pass it to API calls.
const khr_external_memory_capabilities = 1
pub const khr_external_memory_capabilities_spec_version = 1
pub const khr_external_memory_capabilities_extension_name = "VK_KHR_external_memory_capabilities"
pub const luid_size_khr                     = luid_size
pub type ExternalMemoryHandleTypeFlagBitsKHR = ExternalMemoryHandleTypeFlagBits

pub type ExternalMemoryFeatureFlagBitsKHR = ExternalMemoryFeatureFlagBits

pub type ExternalMemoryPropertiesKHR = ExternalMemoryProperties

pub type PhysicalDeviceExternalImageFormatInfoKHR = PhysicalDeviceExternalImageFormatInfo

pub type ExternalImageFormatPropertiesKHR = ExternalImageFormatProperties

pub type PhysicalDeviceExternalBufferInfoKHR = PhysicalDeviceExternalBufferInfo

pub type ExternalBufferPropertiesKHR = ExternalBufferProperties

pub type PhysicalDeviceIDPropertiesKHR = PhysicalDeviceIDProperties

type VkGetPhysicalDeviceExternalBufferPropertiesKHR = fn (     C.PhysicalDevice,     &PhysicalDeviceExternalBufferInfo,     &ExternalBufferProperties) 

pub fn get_physical_device_external_buffer_properties_khr(
    physical_device                                 C.PhysicalDevice,
    p_external_buffer_info                          &PhysicalDeviceExternalBufferInfo,
    p_external_buffer_properties                    &ExternalBufferProperties)  {
      f := VkGetPhysicalDeviceExternalBufferPropertiesKHR((*loader_p).get_sym('vkGetPhysicalDeviceExternalBufferPropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceExternalBufferPropertiesKHR': ${err}")
        return 
    })
    f(
    physical_device,
    p_external_buffer_info,
    p_external_buffer_properties)
}




// VK_KHR_external_memory is a preprocessor guard. Do not pass it to API calls.
const khr_external_memory = 1
pub const khr_external_memory_spec_version  = 1
pub const khr_external_memory_extension_name = "VK_KHR_external_memory"
pub const queue_family_external_khr         = queue_family_external
pub type ExternalMemoryImageCreateInfoKHR = ExternalMemoryImageCreateInfo

pub type ExternalMemoryBufferCreateInfoKHR = ExternalMemoryBufferCreateInfo

pub type ExportMemoryAllocateInfoKHR = ExportMemoryAllocateInfo



// VK_KHR_external_memory_win32 is a preprocessor guard. Do not pass it to API calls.
const khr_external_memory_win32 = 1
pub const khr_external_memory_win32_spec_version = 1
pub const khr_external_memory_win32_extension_name = "VK_KHR_external_memory_win32"
// ImportMemoryWin32HandleInfoKHR extends VkMemoryAllocateInfo
pub struct ImportMemoryWin32HandleInfoKHR {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    handle_type                               ExternalMemoryHandleTypeFlagBits
    handle                                    voidptr
    name                                      string
} 

// ExportMemoryWin32HandleInfoKHR extends VkMemoryAllocateInfo
pub struct ExportMemoryWin32HandleInfoKHR {
mut:
    s_type                            StructureType
    p_next                            voidptr
    p_attributes                      voidptr
    dw_access                         u32
    name                              string
} 

pub struct MemoryWin32HandlePropertiesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    memory_type_bits       u32
} 

pub struct MemoryGetWin32HandleInfoKHR {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    memory                                    C.DeviceMemory
    handle_type                               ExternalMemoryHandleTypeFlagBits
} 

type VkGetMemoryWin32HandleKHR = fn (     C.Device,     &MemoryGetWin32HandleInfoKHR,     &voidptr) Result

pub fn get_memory_win32_handle_khr(
    device                                          C.Device,
    p_get_win32_handle_info                         &MemoryGetWin32HandleInfoKHR,
    p_handle                                        &voidptr) Result {
      f := VkGetMemoryWin32HandleKHR((*loader_p).get_sym('vkGetMemoryWin32HandleKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetMemoryWin32HandleKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_get_win32_handle_info,
    p_handle)
}


type VkGetMemoryWin32HandlePropertiesKHR = fn (     C.Device,     ExternalMemoryHandleTypeFlagBits,     voidptr,     &MemoryWin32HandlePropertiesKHR) Result

pub fn get_memory_win32_handle_properties_khr(
    device                                          C.Device,
    handle_type                                     ExternalMemoryHandleTypeFlagBits,
    handle                                          voidptr,
    p_memory_win32_handle_properties                &MemoryWin32HandlePropertiesKHR) Result {
      f := VkGetMemoryWin32HandlePropertiesKHR((*loader_p).get_sym('vkGetMemoryWin32HandlePropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetMemoryWin32HandlePropertiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    handle_type,
    handle,
    p_memory_win32_handle_properties)
}




// VK_KHR_external_memory_fd is a preprocessor guard. Do not pass it to API calls.
const khr_external_memory_fd = 1
pub const khr_external_memory_fd_spec_version = 1
pub const khr_external_memory_fd_extension_name = "VK_KHR_external_memory_fd"
// ImportMemoryFdInfoKHR extends VkMemoryAllocateInfo
pub struct ImportMemoryFdInfoKHR {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    handle_type                               ExternalMemoryHandleTypeFlagBits
    fd                                        int
} 

pub struct MemoryFdPropertiesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    memory_type_bits       u32
} 

pub struct MemoryGetFdInfoKHR {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    memory                                    C.DeviceMemory
    handle_type                               ExternalMemoryHandleTypeFlagBits
} 

type VkGetMemoryFdKHR = fn (     C.Device,     &MemoryGetFdInfoKHR,     &int) Result

pub fn get_memory_fd_khr(
    device                                          C.Device,
    p_get_fd_info                                   &MemoryGetFdInfoKHR,
    p_fd                                            &int) Result {
      f := VkGetMemoryFdKHR((*loader_p).get_sym('vkGetMemoryFdKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetMemoryFdKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_get_fd_info,
    p_fd)
}


type VkGetMemoryFdPropertiesKHR = fn (     C.Device,     ExternalMemoryHandleTypeFlagBits,     int,     &MemoryFdPropertiesKHR) Result

pub fn get_memory_fd_properties_khr(
    device                                          C.Device,
    handle_type                                     ExternalMemoryHandleTypeFlagBits,
    fd                                              int,
    p_memory_fd_properties                          &MemoryFdPropertiesKHR) Result {
      f := VkGetMemoryFdPropertiesKHR((*loader_p).get_sym('vkGetMemoryFdPropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetMemoryFdPropertiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    handle_type,
    fd,
    p_memory_fd_properties)
}




// VK_KHR_win32_keyed_mutex is a preprocessor guard. Do not pass it to API calls.
const khr_win32_keyed_mutex = 1
pub const khr_win32_keyed_mutex_spec_version = 1
pub const khr_win32_keyed_mutex_extension_name = "VK_KHR_win32_keyed_mutex"
// Win32KeyedMutexAcquireReleaseInfoKHR extends VkSubmitInfo,VkSubmitInfo2
pub struct Win32KeyedMutexAcquireReleaseInfoKHR {
mut:
    s_type                       StructureType
    p_next                       voidptr
    acquire_count                u32
    p_acquire_syncs              &C.DeviceMemory
    p_acquire_keys               &u64
    p_acquire_timeouts           &u32
    release_count                u32
    p_release_syncs              &C.DeviceMemory
    p_release_keys               &u64
} 



// VK_KHR_external_semaphore_capabilities is a preprocessor guard. Do not pass it to API calls.
const khr_external_semaphore_capabilities = 1
pub const khr_external_semaphore_capabilities_spec_version = 1
pub const khr_external_semaphore_capabilities_extension_name = "VK_KHR_external_semaphore_capabilities"
pub type ExternalSemaphoreHandleTypeFlagBitsKHR = ExternalSemaphoreHandleTypeFlagBits

pub type ExternalSemaphoreFeatureFlagBitsKHR = ExternalSemaphoreFeatureFlagBits

pub type PhysicalDeviceExternalSemaphoreInfoKHR = PhysicalDeviceExternalSemaphoreInfo

pub type ExternalSemaphorePropertiesKHR = ExternalSemaphoreProperties

type VkGetPhysicalDeviceExternalSemaphorePropertiesKHR = fn (     C.PhysicalDevice,     &PhysicalDeviceExternalSemaphoreInfo,     &ExternalSemaphoreProperties) 

pub fn get_physical_device_external_semaphore_properties_khr(
    physical_device                                 C.PhysicalDevice,
    p_external_semaphore_info                       &PhysicalDeviceExternalSemaphoreInfo,
    p_external_semaphore_properties                 &ExternalSemaphoreProperties)  {
      f := VkGetPhysicalDeviceExternalSemaphorePropertiesKHR((*loader_p).get_sym('vkGetPhysicalDeviceExternalSemaphorePropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceExternalSemaphorePropertiesKHR': ${err}")
        return 
    })
    f(
    physical_device,
    p_external_semaphore_info,
    p_external_semaphore_properties)
}




// VK_KHR_external_semaphore is a preprocessor guard. Do not pass it to API calls.
const khr_external_semaphore = 1
pub const khr_external_semaphore_spec_version = 1
pub const khr_external_semaphore_extension_name = "VK_KHR_external_semaphore"
pub type SemaphoreImportFlagBitsKHR = SemaphoreImportFlagBits

pub type ExportSemaphoreCreateInfoKHR = ExportSemaphoreCreateInfo



// VK_KHR_external_semaphore_win32 is a preprocessor guard. Do not pass it to API calls.
const khr_external_semaphore_win32 = 1
pub const khr_external_semaphore_win32_spec_version = 1
pub const khr_external_semaphore_win32_extension_name = "VK_KHR_external_semaphore_win32"
pub struct ImportSemaphoreWin32HandleInfoKHR {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    semaphore                                    C.Semaphore
    flags                                        SemaphoreImportFlags
    handle_type                                  ExternalSemaphoreHandleTypeFlagBits
    handle                                       voidptr
    name                                         string
} 

// ExportSemaphoreWin32HandleInfoKHR extends VkSemaphoreCreateInfo
pub struct ExportSemaphoreWin32HandleInfoKHR {
mut:
    s_type                            StructureType
    p_next                            voidptr
    p_attributes                      voidptr
    dw_access                         u32
    name                              string
} 

// D3D12FenceSubmitInfoKHR extends VkSubmitInfo
pub struct D3D12FenceSubmitInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    wait_semaphore_values_count u32
    p_wait_semaphore_values &u64
    signal_semaphore_values_count u32
    p_signal_semaphore_values &u64
} 

pub struct SemaphoreGetWin32HandleInfoKHR {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    semaphore                                    C.Semaphore
    handle_type                                  ExternalSemaphoreHandleTypeFlagBits
} 

type VkImportSemaphoreWin32HandleKHR = fn (     C.Device,     &ImportSemaphoreWin32HandleInfoKHR) Result

pub fn import_semaphore_win32_handle_khr(
    device                                          C.Device,
    p_import_semaphore_win32_handle_info            &ImportSemaphoreWin32HandleInfoKHR) Result {
      f := VkImportSemaphoreWin32HandleKHR((*loader_p).get_sym('vkImportSemaphoreWin32HandleKHR'
    ) or { 
        println("Couldn't load symbol for 'vkImportSemaphoreWin32HandleKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_import_semaphore_win32_handle_info)
}


type VkGetSemaphoreWin32HandleKHR = fn (     C.Device,     &SemaphoreGetWin32HandleInfoKHR,     &voidptr) Result

pub fn get_semaphore_win32_handle_khr(
    device                                          C.Device,
    p_get_win32_handle_info                         &SemaphoreGetWin32HandleInfoKHR,
    p_handle                                        &voidptr) Result {
      f := VkGetSemaphoreWin32HandleKHR((*loader_p).get_sym('vkGetSemaphoreWin32HandleKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetSemaphoreWin32HandleKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_get_win32_handle_info,
    p_handle)
}




// VK_KHR_external_semaphore_fd is a preprocessor guard. Do not pass it to API calls.
const khr_external_semaphore_fd = 1
pub const khr_external_semaphore_fd_spec_version = 1
pub const khr_external_semaphore_fd_extension_name = "VK_KHR_external_semaphore_fd"
pub struct ImportSemaphoreFdInfoKHR {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    semaphore                                    C.Semaphore
    flags                                        SemaphoreImportFlags
    handle_type                                  ExternalSemaphoreHandleTypeFlagBits
    fd                                           int
} 

pub struct SemaphoreGetFdInfoKHR {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    semaphore                                    C.Semaphore
    handle_type                                  ExternalSemaphoreHandleTypeFlagBits
} 

type VkImportSemaphoreFdKHR = fn (     C.Device,     &ImportSemaphoreFdInfoKHR) Result

pub fn import_semaphore_fd_khr(
    device                                          C.Device,
    p_import_semaphore_fd_info                      &ImportSemaphoreFdInfoKHR) Result {
      f := VkImportSemaphoreFdKHR((*loader_p).get_sym('vkImportSemaphoreFdKHR'
    ) or { 
        println("Couldn't load symbol for 'vkImportSemaphoreFdKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_import_semaphore_fd_info)
}


type VkGetSemaphoreFdKHR = fn (     C.Device,     &SemaphoreGetFdInfoKHR,     &int) Result

pub fn get_semaphore_fd_khr(
    device                                          C.Device,
    p_get_fd_info                                   &SemaphoreGetFdInfoKHR,
    p_fd                                            &int) Result {
      f := VkGetSemaphoreFdKHR((*loader_p).get_sym('vkGetSemaphoreFdKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetSemaphoreFdKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_get_fd_info,
    p_fd)
}




// VK_KHR_push_descriptor is a preprocessor guard. Do not pass it to API calls.
const khr_push_descriptor = 1
pub const khr_push_descriptor_spec_version  = 2
pub const khr_push_descriptor_extension_name = "VK_KHR_push_descriptor"
// PhysicalDevicePushDescriptorPropertiesKHR extends VkPhysicalDeviceProperties2
pub struct PhysicalDevicePushDescriptorPropertiesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_push_descriptors   u32
} 

type VkCmdPushDescriptorSetKHR = fn (     C.CommandBuffer,     PipelineBindPoint,     C.PipelineLayout,     u32,     u32,     &WriteDescriptorSet) 

pub fn cmd_push_descriptor_set_khr(
    command_buffer                                  C.CommandBuffer,
    pipeline_bind_point                             PipelineBindPoint,
    layout                                          C.PipelineLayout,
    set                                             u32,
    descriptor_write_count                          u32,
    p_descriptor_writes                             &WriteDescriptorSet)  {
      f := VkCmdPushDescriptorSetKHR((*loader_p).get_sym('vkCmdPushDescriptorSetKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdPushDescriptorSetKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    pipeline_bind_point,
    layout,
    set,
    descriptor_write_count,
    p_descriptor_writes)
}


type VkCmdPushDescriptorSetWithTemplateKHR = fn (     C.CommandBuffer,     C.DescriptorUpdateTemplate,     C.PipelineLayout,     u32,     voidptr) 

pub fn cmd_push_descriptor_set_with_template_khr(
    command_buffer                                  C.CommandBuffer,
    descriptor_update_template                      C.DescriptorUpdateTemplate,
    layout                                          C.PipelineLayout,
    set                                             u32,
    p_data                                          voidptr)  {
      f := VkCmdPushDescriptorSetWithTemplateKHR((*loader_p).get_sym('vkCmdPushDescriptorSetWithTemplateKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdPushDescriptorSetWithTemplateKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    descriptor_update_template,
    layout,
    set,
    p_data)
}




// VK_KHR_shader_float16_int8 is a preprocessor guard. Do not pass it to API calls.
const khr_shader_float16_int8 = 1
pub const khr_shader_float16_int8_spec_version = 1
pub const khr_shader_float16_int8_extension_name = "VK_KHR_shader_float16_int8"
pub type PhysicalDeviceShaderFloat16Int8FeaturesKHR = PhysicalDeviceShaderFloat16Int8Features

pub type PhysicalDeviceFloat16Int8FeaturesKHR = PhysicalDeviceShaderFloat16Int8Features



// VK_KHR_16bit_storage is a preprocessor guard. Do not pass it to API calls.
const khr_16bit_storage = 1
pub const khr_16bit_storage_spec_version    = 1
pub const khr_16bit_storage_extension_name  = "VK_KHR_16bit_storage"
pub type PhysicalDevice16BitStorageFeaturesKHR = PhysicalDevice16BitStorageFeatures



// VK_KHR_incremental_present is a preprocessor guard. Do not pass it to API calls.
const khr_incremental_present = 1
pub const khr_incremental_present_spec_version = 2
pub const khr_incremental_present_extension_name = "VK_KHR_incremental_present"
pub struct RectLayerKHR {
mut:
    offset            Offset2D
    extent            Extent2D
    layer             u32
} 

pub struct PresentRegionKHR {
mut:
    rectangle_count              u32
    p_rectangles                 &RectLayerKHR
} 

// PresentRegionsKHR extends VkPresentInfoKHR
pub struct PresentRegionsKHR {
mut:
    s_type                           StructureType
    p_next                           voidptr
    swapchain_count                  u32
    p_regions                        &PresentRegionKHR
} 



// VK_KHR_descriptor_update_template is a preprocessor guard. Do not pass it to API calls.
const khr_descriptor_update_template = 1
pub const khr_descriptor_update_template_spec_version = 1
pub const khr_descriptor_update_template_extension_name = "VK_KHR_descriptor_update_template"
pub type DescriptorUpdateTemplateTypeKHR = DescriptorUpdateTemplateType

pub type DescriptorUpdateTemplateEntryKHR = DescriptorUpdateTemplateEntry

pub type DescriptorUpdateTemplateCreateInfoKHR = DescriptorUpdateTemplateCreateInfo

type VkCreateDescriptorUpdateTemplateKHR = fn (     C.Device,     &DescriptorUpdateTemplateCreateInfo,     &AllocationCallbacks,     &C.DescriptorUpdateTemplate) Result

pub fn create_descriptor_update_template_khr(
    device                                          C.Device,
    p_create_info                                   &DescriptorUpdateTemplateCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_descriptor_update_template                    &C.DescriptorUpdateTemplate) Result {
      f := VkCreateDescriptorUpdateTemplateKHR((*loader_p).get_sym('vkCreateDescriptorUpdateTemplateKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateDescriptorUpdateTemplateKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_descriptor_update_template)
}


type VkDestroyDescriptorUpdateTemplateKHR = fn (     C.Device,     C.DescriptorUpdateTemplate,     &AllocationCallbacks) 

pub fn destroy_descriptor_update_template_khr(
    device                                          C.Device,
    descriptor_update_template                      C.DescriptorUpdateTemplate,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyDescriptorUpdateTemplateKHR((*loader_p).get_sym('vkDestroyDescriptorUpdateTemplateKHR'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyDescriptorUpdateTemplateKHR': ${err}")
        return 
    })
    f(
    device,
    descriptor_update_template,
    p_allocator)
}


type VkUpdateDescriptorSetWithTemplateKHR = fn (     C.Device,     C.DescriptorSet,     C.DescriptorUpdateTemplate,     voidptr) 

pub fn update_descriptor_set_with_template_khr(
    device                                          C.Device,
    descriptor_set                                  C.DescriptorSet,
    descriptor_update_template                      C.DescriptorUpdateTemplate,
    p_data                                          voidptr)  {
      f := VkUpdateDescriptorSetWithTemplateKHR((*loader_p).get_sym('vkUpdateDescriptorSetWithTemplateKHR'
    ) or { 
        println("Couldn't load symbol for 'vkUpdateDescriptorSetWithTemplateKHR': ${err}")
        return 
    })
    f(
    device,
    descriptor_set,
    descriptor_update_template,
    p_data)
}




// VK_KHR_imageless_framebuffer is a preprocessor guard. Do not pass it to API calls.
const khr_imageless_framebuffer = 1
pub const khr_imageless_framebuffer_spec_version = 1
pub const khr_imageless_framebuffer_extension_name = "VK_KHR_imageless_framebuffer"
pub type PhysicalDeviceImagelessFramebufferFeaturesKHR = PhysicalDeviceImagelessFramebufferFeatures

pub type FramebufferAttachmentsCreateInfoKHR = FramebufferAttachmentsCreateInfo

pub type FramebufferAttachmentImageInfoKHR = FramebufferAttachmentImageInfo

pub type RenderPassAttachmentBeginInfoKHR = RenderPassAttachmentBeginInfo



// VK_KHR_create_renderpass2 is a preprocessor guard. Do not pass it to API calls.
const khr_create_renderpass2 = 1
pub const khr_create_renderpass_2_spec_version = 1
pub const khr_create_renderpass_2_extension_name = "VK_KHR_create_renderpass2"
pub type RenderPassCreateInfo2KHR = RenderPassCreateInfo2

pub type AttachmentDescription2KHR = AttachmentDescription2

pub type AttachmentReference2KHR = AttachmentReference2

pub type SubpassDescription2KHR = SubpassDescription2

pub type SubpassDependency2KHR = SubpassDependency2

pub type SubpassBeginInfoKHR = SubpassBeginInfo

pub type SubpassEndInfoKHR = SubpassEndInfo

type VkCreateRenderPass2KHR = fn (     C.Device,     &RenderPassCreateInfo2,     &AllocationCallbacks,     &C.RenderPass) Result

pub fn create_render_pass2_khr(
    device                                          C.Device,
    p_create_info                                   &RenderPassCreateInfo2,
    p_allocator                                     &AllocationCallbacks,
    p_render_pass                                   &C.RenderPass) Result {
      f := VkCreateRenderPass2KHR((*loader_p).get_sym('vkCreateRenderPass2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateRenderPass2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_render_pass)
}


type VkCmdBeginRenderPass2KHR = fn (     C.CommandBuffer,     &RenderPassBeginInfo,     &SubpassBeginInfo) 

pub fn cmd_begin_render_pass2_khr(
    command_buffer                                  C.CommandBuffer,
    p_render_pass_begin                             &RenderPassBeginInfo,
    p_subpass_begin_info                            &SubpassBeginInfo)  {
      f := VkCmdBeginRenderPass2KHR((*loader_p).get_sym('vkCmdBeginRenderPass2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBeginRenderPass2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_render_pass_begin,
    p_subpass_begin_info)
}


type VkCmdNextSubpass2KHR = fn (     C.CommandBuffer,     &SubpassBeginInfo,     &SubpassEndInfo) 

pub fn cmd_next_subpass2_khr(
    command_buffer                                  C.CommandBuffer,
    p_subpass_begin_info                            &SubpassBeginInfo,
    p_subpass_end_info                              &SubpassEndInfo)  {
      f := VkCmdNextSubpass2KHR((*loader_p).get_sym('vkCmdNextSubpass2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdNextSubpass2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_subpass_begin_info,
    p_subpass_end_info)
}


type VkCmdEndRenderPass2KHR = fn (     C.CommandBuffer,     &SubpassEndInfo) 

pub fn cmd_end_render_pass2_khr(
    command_buffer                                  C.CommandBuffer,
    p_subpass_end_info                              &SubpassEndInfo)  {
      f := VkCmdEndRenderPass2KHR((*loader_p).get_sym('vkCmdEndRenderPass2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEndRenderPass2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_subpass_end_info)
}




// VK_KHR_shared_presentable_image is a preprocessor guard. Do not pass it to API calls.
const khr_shared_presentable_image = 1
pub const khr_shared_presentable_image_spec_version = 1
pub const khr_shared_presentable_image_extension_name = "VK_KHR_shared_presentable_image"
// SharedPresentSurfaceCapabilitiesKHR extends VkSurfaceCapabilities2KHR
pub struct SharedPresentSurfaceCapabilitiesKHR {
mut:
    s_type                   StructureType
    p_next                   voidptr
    shared_present_supported_usage_flags ImageUsageFlags
} 

type VkGetSwapchainStatusKHR = fn (     C.Device,     C.SwapchainKHR) Result

pub fn get_swapchain_status_khr(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR) Result {
      f := VkGetSwapchainStatusKHR((*loader_p).get_sym('vkGetSwapchainStatusKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetSwapchainStatusKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain)
}




// VK_KHR_external_fence_capabilities is a preprocessor guard. Do not pass it to API calls.
const khr_external_fence_capabilities = 1
pub const khr_external_fence_capabilities_spec_version = 1
pub const khr_external_fence_capabilities_extension_name = "VK_KHR_external_fence_capabilities"
pub type ExternalFenceHandleTypeFlagBitsKHR = ExternalFenceHandleTypeFlagBits

pub type ExternalFenceFeatureFlagBitsKHR = ExternalFenceFeatureFlagBits

pub type PhysicalDeviceExternalFenceInfoKHR = PhysicalDeviceExternalFenceInfo

pub type ExternalFencePropertiesKHR = ExternalFenceProperties

type VkGetPhysicalDeviceExternalFencePropertiesKHR = fn (     C.PhysicalDevice,     &PhysicalDeviceExternalFenceInfo,     &ExternalFenceProperties) 

pub fn get_physical_device_external_fence_properties_khr(
    physical_device                                 C.PhysicalDevice,
    p_external_fence_info                           &PhysicalDeviceExternalFenceInfo,
    p_external_fence_properties                     &ExternalFenceProperties)  {
      f := VkGetPhysicalDeviceExternalFencePropertiesKHR((*loader_p).get_sym('vkGetPhysicalDeviceExternalFencePropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceExternalFencePropertiesKHR': ${err}")
        return 
    })
    f(
    physical_device,
    p_external_fence_info,
    p_external_fence_properties)
}




// VK_KHR_external_fence is a preprocessor guard. Do not pass it to API calls.
const khr_external_fence = 1
pub const khr_external_fence_spec_version   = 1
pub const khr_external_fence_extension_name = "VK_KHR_external_fence"
pub type FenceImportFlagBitsKHR = FenceImportFlagBits

pub type ExportFenceCreateInfoKHR = ExportFenceCreateInfo



// VK_KHR_external_fence_win32 is a preprocessor guard. Do not pass it to API calls.
const khr_external_fence_win32 = 1
pub const khr_external_fence_win32_spec_version = 1
pub const khr_external_fence_win32_extension_name = "VK_KHR_external_fence_win32"
pub struct ImportFenceWin32HandleInfoKHR {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    fence                                    C.Fence
    flags                                    FenceImportFlags
    handle_type                              ExternalFenceHandleTypeFlagBits
    handle                                   voidptr
    name                                     string
} 

// ExportFenceWin32HandleInfoKHR extends VkFenceCreateInfo
pub struct ExportFenceWin32HandleInfoKHR {
mut:
    s_type                            StructureType
    p_next                            voidptr
    p_attributes                      voidptr
    dw_access                         u32
    name                              string
} 

pub struct FenceGetWin32HandleInfoKHR {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    fence                                    C.Fence
    handle_type                              ExternalFenceHandleTypeFlagBits
} 

type VkImportFenceWin32HandleKHR = fn (     C.Device,     &ImportFenceWin32HandleInfoKHR) Result

pub fn import_fence_win32_handle_khr(
    device                                          C.Device,
    p_import_fence_win32_handle_info                &ImportFenceWin32HandleInfoKHR) Result {
      f := VkImportFenceWin32HandleKHR((*loader_p).get_sym('vkImportFenceWin32HandleKHR'
    ) or { 
        println("Couldn't load symbol for 'vkImportFenceWin32HandleKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_import_fence_win32_handle_info)
}


type VkGetFenceWin32HandleKHR = fn (     C.Device,     &FenceGetWin32HandleInfoKHR,     &voidptr) Result

pub fn get_fence_win32_handle_khr(
    device                                          C.Device,
    p_get_win32_handle_info                         &FenceGetWin32HandleInfoKHR,
    p_handle                                        &voidptr) Result {
      f := VkGetFenceWin32HandleKHR((*loader_p).get_sym('vkGetFenceWin32HandleKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetFenceWin32HandleKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_get_win32_handle_info,
    p_handle)
}




// VK_KHR_external_fence_fd is a preprocessor guard. Do not pass it to API calls.
const khr_external_fence_fd = 1
pub const khr_external_fence_fd_spec_version = 1
pub const khr_external_fence_fd_extension_name = "VK_KHR_external_fence_fd"
pub struct ImportFenceFdInfoKHR {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    fence                                    C.Fence
    flags                                    FenceImportFlags
    handle_type                              ExternalFenceHandleTypeFlagBits
    fd                                       int
} 

pub struct FenceGetFdInfoKHR {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    fence                                    C.Fence
    handle_type                              ExternalFenceHandleTypeFlagBits
} 

type VkImportFenceFdKHR = fn (     C.Device,     &ImportFenceFdInfoKHR) Result

pub fn import_fence_fd_khr(
    device                                          C.Device,
    p_import_fence_fd_info                          &ImportFenceFdInfoKHR) Result {
      f := VkImportFenceFdKHR((*loader_p).get_sym('vkImportFenceFdKHR'
    ) or { 
        println("Couldn't load symbol for 'vkImportFenceFdKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_import_fence_fd_info)
}


type VkGetFenceFdKHR = fn (     C.Device,     &FenceGetFdInfoKHR,     &int) Result

pub fn get_fence_fd_khr(
    device                                          C.Device,
    p_get_fd_info                                   &FenceGetFdInfoKHR,
    p_fd                                            &int) Result {
      f := VkGetFenceFdKHR((*loader_p).get_sym('vkGetFenceFdKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetFenceFdKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_get_fd_info,
    p_fd)
}




// VK_KHR_performance_query is a preprocessor guard. Do not pass it to API calls.
const khr_performance_query = 1
pub const khr_performance_query_spec_version = 1
pub const khr_performance_query_extension_name = "VK_KHR_performance_query"

pub enum PerformanceCounterUnitKHR {
    performance_counter_unit_generic_khr = int(0)
    performance_counter_unit_percentage_khr = int(1)
    performance_counter_unit_nanoseconds_khr = int(2)
    performance_counter_unit_bytes_khr = int(3)
    performance_counter_unit_bytes_per_second_khr = int(4)
    performance_counter_unit_kelvin_khr = int(5)
    performance_counter_unit_watts_khr = int(6)
    performance_counter_unit_volts_khr = int(7)
    performance_counter_unit_amps_khr = int(8)
    performance_counter_unit_hertz_khr = int(9)
    performance_counter_unit_cycles_khr = int(10)
    performance_counter_unit_max_enum_khr = int(0x7FFFFFFF)
}


pub enum PerformanceCounterScopeKHR {
    performance_counter_scope_command_buffer_khr = int(0)
    performance_counter_scope_render_pass_khr = int(1)
    performance_counter_scope_command_khr = int(2)
    performance_counter_scope_max_enum_khr = int(0x7FFFFFFF)
}


pub enum PerformanceCounterStorageKHR {
    performance_counter_storage_int32_khr = int(0)
    performance_counter_storage_int64_khr = int(1)
    performance_counter_storage_uint32_khr = int(2)
    performance_counter_storage_uint64_khr = int(3)
    performance_counter_storage_float32_khr = int(4)
    performance_counter_storage_float64_khr = int(5)
    performance_counter_storage_max_enum_khr = int(0x7FFFFFFF)
}


pub enum PerformanceCounterDescriptionFlagBitsKHR {
    performance_counter_description_performance_impacting_bit_khr = int(0x00000001)
    performance_counter_description_concurrently_impacted_bit_khr = int(0x00000002)
    performance_counter_description_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type PerformanceCounterDescriptionFlagsKHR = u32

pub enum AcquireProfilingLockFlagBitsKHR {
    acquire_profiling_lock_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type AcquireProfilingLockFlagsKHR = u32
// PhysicalDevicePerformanceQueryFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePerformanceQueryFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    performance_counter_query_pools Bool32
    performance_counter_multiple_query_pools Bool32
} 

// PhysicalDevicePerformanceQueryPropertiesKHR extends VkPhysicalDeviceProperties2
pub struct PhysicalDevicePerformanceQueryPropertiesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    allow_command_buffer_query_copies Bool32
} 

pub struct PerformanceCounterKHR {
mut:
    s_type                                StructureType
    p_next                                voidptr
    unit                                  PerformanceCounterUnitKHR
    scope                                 PerformanceCounterScopeKHR
    storage                               PerformanceCounterStorageKHR
    uuid                                  []u8
} 

pub struct PerformanceCounterDescriptionKHR {
mut:
    s_type                                         StructureType
    p_next                                         voidptr
    flags                                          PerformanceCounterDescriptionFlagsKHR
    name                                           []char
    category                                       []char
    description                                    []char
} 

// QueryPoolPerformanceCreateInfoKHR extends VkQueryPoolCreateInfo
pub struct QueryPoolPerformanceCreateInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    queue_family_index     u32
    counter_index_count    u32
    p_counter_indices      &u32
} 

pub union PerformanceCounterResultKHR {
mut:
    int32           i32
    int64           i64
    uint32          u32
    uint64          u64
    float32         f32
    float64         f64
} 

pub struct AcquireProfilingLockInfoKHR {
mut:
    s_type                                StructureType
    p_next                                voidptr
    flags                                 AcquireProfilingLockFlagsKHR
    timeout                               u64
} 

// PerformanceQuerySubmitInfoKHR extends VkSubmitInfo,VkSubmitInfo2
pub struct PerformanceQuerySubmitInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    counter_pass_index     u32
} 

type VkEnumeratePhysicalDeviceQueueFamilyPerformanceQueryCountersKHR = fn (     C.PhysicalDevice,     u32,     &u32,     &PerformanceCounterKHR,     &PerformanceCounterDescriptionKHR) Result

pub fn enumerate_physical_device_queue_family_performance_query_counters_khr(
    physical_device                                 C.PhysicalDevice,
    queue_family_index                              u32,
    p_counter_count                                 &u32,
    p_counters                                      &PerformanceCounterKHR,
    p_counter_descriptions                          &PerformanceCounterDescriptionKHR) Result {
      f := VkEnumeratePhysicalDeviceQueueFamilyPerformanceQueryCountersKHR((*loader_p).get_sym('vkEnumeratePhysicalDeviceQueueFamilyPerformanceQueryCountersKHR'
    ) or { 
        println("Couldn't load symbol for 'vkEnumeratePhysicalDeviceQueueFamilyPerformanceQueryCountersKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    queue_family_index,
    p_counter_count,
    p_counters,
    p_counter_descriptions)
}


type VkGetPhysicalDeviceQueueFamilyPerformanceQueryPassesKHR = fn (     C.PhysicalDevice,     &QueryPoolPerformanceCreateInfoKHR,     &u32) 

pub fn get_physical_device_queue_family_performance_query_passes_khr(
    physical_device                                 C.PhysicalDevice,
    p_performance_query_create_info                 &QueryPoolPerformanceCreateInfoKHR,
    p_num_passes                                    &u32)  {
      f := VkGetPhysicalDeviceQueueFamilyPerformanceQueryPassesKHR((*loader_p).get_sym('vkGetPhysicalDeviceQueueFamilyPerformanceQueryPassesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceQueueFamilyPerformanceQueryPassesKHR': ${err}")
        return 
    })
    f(
    physical_device,
    p_performance_query_create_info,
    p_num_passes)
}


type VkAcquireProfilingLockKHR = fn (     C.Device,     &AcquireProfilingLockInfoKHR) Result

pub fn acquire_profiling_lock_khr(
    device                                          C.Device,
    p_info                                          &AcquireProfilingLockInfoKHR) Result {
      f := VkAcquireProfilingLockKHR((*loader_p).get_sym('vkAcquireProfilingLockKHR'
    ) or { 
        println("Couldn't load symbol for 'vkAcquireProfilingLockKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_info)
}


type VkReleaseProfilingLockKHR = fn (     C.Device) 

pub fn release_profiling_lock_khr(
    device                                          C.Device)  {
      f := VkReleaseProfilingLockKHR((*loader_p).get_sym('vkReleaseProfilingLockKHR'
    ) or { 
        println("Couldn't load symbol for 'vkReleaseProfilingLockKHR': ${err}")
        return 
    })
    f(
    device)
}




// VK_KHR_maintenance2 is a preprocessor guard. Do not pass it to API calls.
const khr_maintenance2 = 1
pub const khr_maintenance_2_spec_version    = 1
pub const khr_maintenance_2_extension_name  = "VK_KHR_maintenance2"
pub const khr_maintenance2_spec_version     = khr_maintenance_2_spec_version
pub const khr_maintenance2_extension_name   = khr_maintenance_2_extension_name
pub type PointClippingBehaviorKHR = PointClippingBehavior

pub type TessellationDomainOriginKHR = TessellationDomainOrigin

pub type PhysicalDevicePointClippingPropertiesKHR = PhysicalDevicePointClippingProperties

pub type RenderPassInputAttachmentAspectCreateInfoKHR = RenderPassInputAttachmentAspectCreateInfo

pub type InputAttachmentAspectReferenceKHR = InputAttachmentAspectReference

pub type ImageViewUsageCreateInfoKHR = ImageViewUsageCreateInfo

pub type PipelineTessellationDomainOriginStateCreateInfoKHR = PipelineTessellationDomainOriginStateCreateInfo



// VK_KHR_get_surface_capabilities2 is a preprocessor guard. Do not pass it to API calls.
const khr_get_surface_capabilities2 = 1
pub const khr_get_surface_capabilities_2_spec_version = 1
pub const khr_get_surface_capabilities_2_extension_name = "VK_KHR_get_surface_capabilities2"
pub struct PhysicalDeviceSurfaceInfo2KHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    surface                C.SurfaceKHR
} 

pub struct SurfaceCapabilities2KHR {
mut:
    s_type                          StructureType
    p_next                          voidptr
    surface_capabilities            SurfaceCapabilitiesKHR
} 

pub struct SurfaceFormat2KHR {
mut:
    s_type                    StructureType
    p_next                    voidptr
    surface_format            SurfaceFormatKHR
} 

type VkGetPhysicalDeviceSurfaceCapabilities2KHR = fn (     C.PhysicalDevice,     &PhysicalDeviceSurfaceInfo2KHR,     &SurfaceCapabilities2KHR) Result

pub fn get_physical_device_surface_capabilities2_khr(
    physical_device                                 C.PhysicalDevice,
    p_surface_info                                  &PhysicalDeviceSurfaceInfo2KHR,
    p_surface_capabilities                          &SurfaceCapabilities2KHR) Result {
      f := VkGetPhysicalDeviceSurfaceCapabilities2KHR((*loader_p).get_sym('vkGetPhysicalDeviceSurfaceCapabilities2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSurfaceCapabilities2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_surface_info,
    p_surface_capabilities)
}


type VkGetPhysicalDeviceSurfaceFormats2KHR = fn (     C.PhysicalDevice,     &PhysicalDeviceSurfaceInfo2KHR,     &u32,     &SurfaceFormat2KHR) Result

pub fn get_physical_device_surface_formats2_khr(
    physical_device                                 C.PhysicalDevice,
    p_surface_info                                  &PhysicalDeviceSurfaceInfo2KHR,
    p_surface_format_count                          &u32,
    p_surface_formats                               &SurfaceFormat2KHR) Result {
      f := VkGetPhysicalDeviceSurfaceFormats2KHR((*loader_p).get_sym('vkGetPhysicalDeviceSurfaceFormats2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSurfaceFormats2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_surface_info,
    p_surface_format_count,
    p_surface_formats)
}




// VK_KHR_variable_pointers is a preprocessor guard. Do not pass it to API calls.
const khr_variable_pointers = 1
pub const khr_variable_pointers_spec_version = 1
pub const khr_variable_pointers_extension_name = "VK_KHR_variable_pointers"
pub type PhysicalDeviceVariablePointerFeaturesKHR = PhysicalDeviceVariablePointersFeatures

pub type PhysicalDeviceVariablePointersFeaturesKHR = PhysicalDeviceVariablePointersFeatures



// VK_KHR_get_display_properties2 is a preprocessor guard. Do not pass it to API calls.
const khr_get_display_properties2 = 1
pub const khr_get_display_properties_2_spec_version = 1
pub const khr_get_display_properties_2_extension_name = "VK_KHR_get_display_properties2"
pub struct DisplayProperties2KHR {
mut:
    s_type                        StructureType
    p_next                        voidptr
    display_properties            DisplayPropertiesKHR
} 

pub struct DisplayPlaneProperties2KHR {
mut:
    s_type                             StructureType
    p_next                             voidptr
    display_plane_properties           DisplayPlanePropertiesKHR
} 

pub struct DisplayModeProperties2KHR {
mut:
    s_type                            StructureType
    p_next                            voidptr
    display_mode_properties           DisplayModePropertiesKHR
} 

pub struct DisplayPlaneInfo2KHR {
mut:
    s_type                  StructureType
    p_next                  voidptr
    mode                    C.DisplayModeKHR
    plane_index             u32
} 

pub struct DisplayPlaneCapabilities2KHR {
mut:
    s_type                               StructureType
    p_next                               voidptr
    capabilities                         DisplayPlaneCapabilitiesKHR
} 

type VkGetPhysicalDeviceDisplayProperties2KHR = fn (     C.PhysicalDevice,     &u32,     &DisplayProperties2KHR) Result

pub fn get_physical_device_display_properties2_khr(
    physical_device                                 C.PhysicalDevice,
    p_property_count                                &u32,
    p_properties                                    &DisplayProperties2KHR) Result {
      f := VkGetPhysicalDeviceDisplayProperties2KHR((*loader_p).get_sym('vkGetPhysicalDeviceDisplayProperties2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceDisplayProperties2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_property_count,
    p_properties)
}


type VkGetPhysicalDeviceDisplayPlaneProperties2KHR = fn (     C.PhysicalDevice,     &u32,     &DisplayPlaneProperties2KHR) Result

pub fn get_physical_device_display_plane_properties2_khr(
    physical_device                                 C.PhysicalDevice,
    p_property_count                                &u32,
    p_properties                                    &DisplayPlaneProperties2KHR) Result {
      f := VkGetPhysicalDeviceDisplayPlaneProperties2KHR((*loader_p).get_sym('vkGetPhysicalDeviceDisplayPlaneProperties2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceDisplayPlaneProperties2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_property_count,
    p_properties)
}


type VkGetDisplayModeProperties2KHR = fn (     C.PhysicalDevice,     C.DisplayKHR,     &u32,     &DisplayModeProperties2KHR) Result

pub fn get_display_mode_properties2_khr(
    physical_device                                 C.PhysicalDevice,
    display                                         C.DisplayKHR,
    p_property_count                                &u32,
    p_properties                                    &DisplayModeProperties2KHR) Result {
      f := VkGetDisplayModeProperties2KHR((*loader_p).get_sym('vkGetDisplayModeProperties2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDisplayModeProperties2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    display,
    p_property_count,
    p_properties)
}


type VkGetDisplayPlaneCapabilities2KHR = fn (     C.PhysicalDevice,     &DisplayPlaneInfo2KHR,     &DisplayPlaneCapabilities2KHR) Result

pub fn get_display_plane_capabilities2_khr(
    physical_device                                 C.PhysicalDevice,
    p_display_plane_info                            &DisplayPlaneInfo2KHR,
    p_capabilities                                  &DisplayPlaneCapabilities2KHR) Result {
      f := VkGetDisplayPlaneCapabilities2KHR((*loader_p).get_sym('vkGetDisplayPlaneCapabilities2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDisplayPlaneCapabilities2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_display_plane_info,
    p_capabilities)
}




// VK_KHR_dedicated_allocation is a preprocessor guard. Do not pass it to API calls.
const khr_dedicated_allocation = 1
pub const khr_dedicated_allocation_spec_version = 3
pub const khr_dedicated_allocation_extension_name = "VK_KHR_dedicated_allocation"
pub type MemoryDedicatedRequirementsKHR = MemoryDedicatedRequirements

pub type MemoryDedicatedAllocateInfoKHR = MemoryDedicatedAllocateInfo



// VK_KHR_storage_buffer_storage_class is a preprocessor guard. Do not pass it to API calls.
const khr_storage_buffer_storage_class = 1
pub const khr_storage_buffer_storage_class_spec_version = 1
pub const khr_storage_buffer_storage_class_extension_name = "VK_KHR_storage_buffer_storage_class"


// VK_KHR_relaxed_block_layout is a preprocessor guard. Do not pass it to API calls.
const khr_relaxed_block_layout = 1
pub const khr_relaxed_block_layout_spec_version = 1
pub const khr_relaxed_block_layout_extension_name = "VK_KHR_relaxed_block_layout"


// VK_KHR_get_memory_requirements2 is a preprocessor guard. Do not pass it to API calls.
const khr_get_memory_requirements2 = 1
pub const khr_get_memory_requirements_2_spec_version = 1
pub const khr_get_memory_requirements_2_extension_name = "VK_KHR_get_memory_requirements2"
pub type BufferMemoryRequirementsInfo2KHR = BufferMemoryRequirementsInfo2

pub type ImageMemoryRequirementsInfo2KHR = ImageMemoryRequirementsInfo2

pub type ImageSparseMemoryRequirementsInfo2KHR = ImageSparseMemoryRequirementsInfo2

pub type MemoryRequirements2KHR = MemoryRequirements2

pub type SparseImageMemoryRequirements2KHR = SparseImageMemoryRequirements2

type VkGetImageMemoryRequirements2KHR = fn (     C.Device,     &ImageMemoryRequirementsInfo2,     &MemoryRequirements2) 

pub fn get_image_memory_requirements2_khr(
    device                                          C.Device,
    p_info                                          &ImageMemoryRequirementsInfo2,
    p_memory_requirements                           &MemoryRequirements2)  {
      f := VkGetImageMemoryRequirements2KHR((*loader_p).get_sym('vkGetImageMemoryRequirements2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageMemoryRequirements2KHR': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_memory_requirements)
}


type VkGetBufferMemoryRequirements2KHR = fn (     C.Device,     &BufferMemoryRequirementsInfo2,     &MemoryRequirements2) 

pub fn get_buffer_memory_requirements2_khr(
    device                                          C.Device,
    p_info                                          &BufferMemoryRequirementsInfo2,
    p_memory_requirements                           &MemoryRequirements2)  {
      f := VkGetBufferMemoryRequirements2KHR((*loader_p).get_sym('vkGetBufferMemoryRequirements2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetBufferMemoryRequirements2KHR': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_memory_requirements)
}


type VkGetImageSparseMemoryRequirements2KHR = fn (     C.Device,     &ImageSparseMemoryRequirementsInfo2,     &u32,     &SparseImageMemoryRequirements2) 

pub fn get_image_sparse_memory_requirements2_khr(
    device                                          C.Device,
    p_info                                          &ImageSparseMemoryRequirementsInfo2,
    p_sparse_memory_requirement_count               &u32,
    p_sparse_memory_requirements                    &SparseImageMemoryRequirements2)  {
      f := VkGetImageSparseMemoryRequirements2KHR((*loader_p).get_sym('vkGetImageSparseMemoryRequirements2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageSparseMemoryRequirements2KHR': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_sparse_memory_requirement_count,
    p_sparse_memory_requirements)
}




// VK_KHR_image_format_list is a preprocessor guard. Do not pass it to API calls.
const khr_image_format_list = 1
pub const khr_image_format_list_spec_version = 1
pub const khr_image_format_list_extension_name = "VK_KHR_image_format_list"
pub type ImageFormatListCreateInfoKHR = ImageFormatListCreateInfo



// VK_KHR_sampler_ycbcr_conversion is a preprocessor guard. Do not pass it to API calls.
const khr_sampler_ycbcr_conversion = 1
pub const khr_sampler_ycbcr_conversion_spec_version = 14
pub const khr_sampler_ycbcr_conversion_extension_name = "VK_KHR_sampler_ycbcr_conversion"
pub type SamplerYcbcrModelConversionKHR = SamplerYcbcrModelConversion

pub type SamplerYcbcrRangeKHR = SamplerYcbcrRange

pub type ChromaLocationKHR = ChromaLocation

pub type SamplerYcbcrConversionCreateInfoKHR = SamplerYcbcrConversionCreateInfo

pub type SamplerYcbcrConversionInfoKHR = SamplerYcbcrConversionInfo

pub type BindImagePlaneMemoryInfoKHR = BindImagePlaneMemoryInfo

pub type ImagePlaneMemoryRequirementsInfoKHR = ImagePlaneMemoryRequirementsInfo

pub type PhysicalDeviceSamplerYcbcrConversionFeaturesKHR = PhysicalDeviceSamplerYcbcrConversionFeatures

pub type SamplerYcbcrConversionImageFormatPropertiesKHR = SamplerYcbcrConversionImageFormatProperties

type VkCreateSamplerYcbcrConversionKHR = fn (     C.Device,     &SamplerYcbcrConversionCreateInfo,     &AllocationCallbacks,     &C.SamplerYcbcrConversion) Result

pub fn create_sampler_ycbcr_conversion_khr(
    device                                          C.Device,
    p_create_info                                   &SamplerYcbcrConversionCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_ycbcr_conversion                              &C.SamplerYcbcrConversion) Result {
      f := VkCreateSamplerYcbcrConversionKHR((*loader_p).get_sym('vkCreateSamplerYcbcrConversionKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateSamplerYcbcrConversionKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_ycbcr_conversion)
}


type VkDestroySamplerYcbcrConversionKHR = fn (     C.Device,     C.SamplerYcbcrConversion,     &AllocationCallbacks) 

pub fn destroy_sampler_ycbcr_conversion_khr(
    device                                          C.Device,
    ycbcr_conversion                                C.SamplerYcbcrConversion,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroySamplerYcbcrConversionKHR((*loader_p).get_sym('vkDestroySamplerYcbcrConversionKHR'
    ) or { 
        println("Couldn't load symbol for 'vkDestroySamplerYcbcrConversionKHR': ${err}")
        return 
    })
    f(
    device,
    ycbcr_conversion,
    p_allocator)
}




// VK_KHR_bind_memory2 is a preprocessor guard. Do not pass it to API calls.
const khr_bind_memory2 = 1
pub const khr_bind_memory_2_spec_version    = 1
pub const khr_bind_memory_2_extension_name  = "VK_KHR_bind_memory2"
pub type BindBufferMemoryInfoKHR = BindBufferMemoryInfo

pub type BindImageMemoryInfoKHR = BindImageMemoryInfo

type VkBindBufferMemory2KHR = fn (     C.Device,     u32,     &BindBufferMemoryInfo) Result

pub fn bind_buffer_memory2_khr(
    device                                          C.Device,
    bind_info_count                                 u32,
    p_bind_infos                                    &BindBufferMemoryInfo) Result {
      f := VkBindBufferMemory2KHR((*loader_p).get_sym('vkBindBufferMemory2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkBindBufferMemory2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    bind_info_count,
    p_bind_infos)
}


type VkBindImageMemory2KHR = fn (     C.Device,     u32,     &BindImageMemoryInfo) Result

pub fn bind_image_memory2_khr(
    device                                          C.Device,
    bind_info_count                                 u32,
    p_bind_infos                                    &BindImageMemoryInfo) Result {
      f := VkBindImageMemory2KHR((*loader_p).get_sym('vkBindImageMemory2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkBindImageMemory2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    bind_info_count,
    p_bind_infos)
}




// VK_KHR_portability_subset is a preprocessor guard. Do not pass it to API calls.
const khr_portability_subset = 1
pub const khr_portability_subset_spec_version = 1
pub const khr_portability_subset_extension_name = "VK_KHR_portability_subset"
// PhysicalDevicePortabilitySubsetFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePortabilitySubsetFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    constant_alpha_color_blend_factors Bool32
    events                 Bool32
    image_view_format_reinterpretation Bool32
    image_view_format_swizzle Bool32
    image_view2_d_on3_d_image Bool32
    multisample_array_image Bool32
    mutable_comparison_samplers Bool32
    point_polygons         Bool32
    sampler_mip_lod_bias   Bool32
    separate_stencil_mask_ref Bool32
    shader_sample_rate_interpolation_functions Bool32
    tessellation_isolines  Bool32
    tessellation_point_mode Bool32
    triangle_fans          Bool32
    vertex_attribute_access_beyond_stride Bool32
} 

// PhysicalDevicePortabilitySubsetPropertiesKHR extends VkPhysicalDeviceProperties2
pub struct PhysicalDevicePortabilitySubsetPropertiesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    min_vertex_input_binding_stride_alignment u32
} 



// VK_KHR_maintenance3 is a preprocessor guard. Do not pass it to API calls.
const khr_maintenance3 = 1
pub const khr_maintenance_3_spec_version    = 1
pub const khr_maintenance_3_extension_name  = "VK_KHR_maintenance3"
pub const khr_maintenance3_spec_version     = khr_maintenance_3_spec_version
pub const khr_maintenance3_extension_name   = khr_maintenance_3_extension_name
pub type PhysicalDeviceMaintenance3PropertiesKHR = PhysicalDeviceMaintenance3Properties

pub type DescriptorSetLayoutSupportKHR = DescriptorSetLayoutSupport

type VkGetDescriptorSetLayoutSupportKHR = fn (     C.Device,     &DescriptorSetLayoutCreateInfo,     &DescriptorSetLayoutSupport) 

pub fn get_descriptor_set_layout_support_khr(
    device                                          C.Device,
    p_create_info                                   &DescriptorSetLayoutCreateInfo,
    p_support                                       &DescriptorSetLayoutSupport)  {
      f := VkGetDescriptorSetLayoutSupportKHR((*loader_p).get_sym('vkGetDescriptorSetLayoutSupportKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDescriptorSetLayoutSupportKHR': ${err}")
        return 
    })
    f(
    device,
    p_create_info,
    p_support)
}




// VK_KHR_draw_indirect_count is a preprocessor guard. Do not pass it to API calls.
const khr_draw_indirect_count = 1
pub const khr_draw_indirect_count_spec_version = 1
pub const khr_draw_indirect_count_extension_name = "VK_KHR_draw_indirect_count"
type VkCmdDrawIndirectCountKHR = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_indirect_count_khr(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    count_buffer                                    C.Buffer,
    count_buffer_offset                             DeviceSize,
    max_draw_count                                  u32,
    stride                                          u32)  {
      f := VkCmdDrawIndirectCountKHR((*loader_p).get_sym('vkCmdDrawIndirectCountKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawIndirectCountKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    count_buffer,
    count_buffer_offset,
    max_draw_count,
    stride)
}


type VkCmdDrawIndexedIndirectCountKHR = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_indexed_indirect_count_khr(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    count_buffer                                    C.Buffer,
    count_buffer_offset                             DeviceSize,
    max_draw_count                                  u32,
    stride                                          u32)  {
      f := VkCmdDrawIndexedIndirectCountKHR((*loader_p).get_sym('vkCmdDrawIndexedIndirectCountKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawIndexedIndirectCountKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    count_buffer,
    count_buffer_offset,
    max_draw_count,
    stride)
}




// VK_KHR_shader_subgroup_extended_types is a preprocessor guard. Do not pass it to API calls.
const khr_shader_subgroup_extended_types = 1
pub const khr_shader_subgroup_extended_types_spec_version = 1
pub const khr_shader_subgroup_extended_types_extension_name = "VK_KHR_shader_subgroup_extended_types"
pub type PhysicalDeviceShaderSubgroupExtendedTypesFeaturesKHR = PhysicalDeviceShaderSubgroupExtendedTypesFeatures



// VK_KHR_8bit_storage is a preprocessor guard. Do not pass it to API calls.
const khr_8bit_storage = 1
pub const khr_8bit_storage_spec_version     = 1
pub const khr_8bit_storage_extension_name   = "VK_KHR_8bit_storage"
pub type PhysicalDevice8BitStorageFeaturesKHR = PhysicalDevice8BitStorageFeatures



// VK_KHR_shader_atomic_int64 is a preprocessor guard. Do not pass it to API calls.
const khr_shader_atomic_int64 = 1
pub const khr_shader_atomic_int64_spec_version = 1
pub const khr_shader_atomic_int64_extension_name = "VK_KHR_shader_atomic_int64"
pub type PhysicalDeviceShaderAtomicInt64FeaturesKHR = PhysicalDeviceShaderAtomicInt64Features



// VK_KHR_shader_clock is a preprocessor guard. Do not pass it to API calls.
const khr_shader_clock = 1
pub const khr_shader_clock_spec_version     = 1
pub const khr_shader_clock_extension_name   = "VK_KHR_shader_clock"
// PhysicalDeviceShaderClockFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderClockFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_subgroup_clock  Bool32
    shader_device_clock    Bool32
} 



// VK_KHR_video_decode_h265 is a preprocessor guard. Do not pass it to API calls.
const khr_video_decode_h265 = 1
pub const khr_video_decode_h265_spec_version = 7
pub const khr_video_decode_h265_extension_name = "VK_KHR_video_decode_h265"
// VideoDecodeH265ProfileInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub struct VideoDecodeH265ProfileInfoKHR {
mut:
    s_type                        StructureType
    p_next                        voidptr
    std_profile_idc               C.StdVideoH265ProfileIdc
} 

// VideoDecodeH265CapabilitiesKHR extends VkVideoCapabilitiesKHR
pub struct VideoDecodeH265CapabilitiesKHR {
mut:
    s_type                      StructureType
    p_next                      voidptr
    max_level_idc               u32
} 

// VideoDecodeH265SessionParametersAddInfoKHR extends VkVideoSessionParametersUpdateInfoKHR
pub struct VideoDecodeH265SessionParametersAddInfoKHR {
mut:
    s_type                                         StructureType
    p_next                                         voidptr
    std_vps_count                                  u32
    p_std_vp_ss                                    &C.StdVideoH265VideoParameterSet
    std_sps_count                                  u32
    p_std_sp_ss                                    &C.StdVideoH265SequenceParameterSet
    std_pps_count                                  u32
    p_std_pp_ss                                    &C.StdVideoH265PictureParameterSet
} 

// VideoDecodeH265SessionParametersCreateInfoKHR extends VkVideoSessionParametersCreateInfoKHR
pub struct VideoDecodeH265SessionParametersCreateInfoKHR {
mut:
    s_type                                                     StructureType
    p_next                                                     voidptr
    max_std_vps_count                                          u32
    max_std_sps_count                                          u32
    max_std_pps_count                                          u32
    p_parameters_add_info                                      &VideoDecodeH265SessionParametersAddInfoKHR
} 

// VideoDecodeH265PictureInfoKHR extends VkVideoDecodeInfoKHR
pub struct VideoDecodeH265PictureInfoKHR {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    p_std_picture_info                          &C.StdVideoDecodeH265PictureInfo
    slice_segment_count                         u32
    p_slice_segment_offsets                     &u32
} 

// VideoDecodeH265DpbSlotInfoKHR extends VkVideoReferenceSlotInfoKHR
pub struct VideoDecodeH265DpbSlotInfoKHR {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    p_std_reference_info                          &C.StdVideoDecodeH265ReferenceInfo
} 



// VK_KHR_global_priority is a preprocessor guard. Do not pass it to API calls.
const khr_global_priority = 1
pub const max_global_priority_size_khr      = u32(16)
pub const khr_global_priority_spec_version  = 1
pub const khr_global_priority_extension_name = "VK_KHR_global_priority"

pub enum QueueGlobalPriorityKHR {
    queue_global_priority_low_khr = int(128)
    queue_global_priority_medium_khr = int(256)
    queue_global_priority_high_khr = int(512)
    queue_global_priority_realtime_khr = int(1024)
    queue_global_priority_max_enum_khr = int(0x7FFFFFFF)
}

// DeviceQueueGlobalPriorityCreateInfoKHR extends VkDeviceQueueCreateInfo
pub struct DeviceQueueGlobalPriorityCreateInfoKHR {
mut:
    s_type                          StructureType
    p_next                          voidptr
    global_priority                 QueueGlobalPriorityKHR
} 

// PhysicalDeviceGlobalPriorityQueryFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceGlobalPriorityQueryFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    global_priority_query  Bool32
} 

// QueueFamilyGlobalPriorityPropertiesKHR extends VkQueueFamilyProperties2
pub struct QueueFamilyGlobalPriorityPropertiesKHR {
mut:
    s_type                          StructureType
    p_next                          voidptr
    priority_count                  u32
    priorities                      []QueueGlobalPriorityKHR
} 



// VK_KHR_driver_properties is a preprocessor guard. Do not pass it to API calls.
const khr_driver_properties = 1
pub const khr_driver_properties_spec_version = 1
pub const khr_driver_properties_extension_name = "VK_KHR_driver_properties"
pub const max_driver_name_size_khr          = max_driver_name_size
pub const max_driver_info_size_khr          = max_driver_info_size
pub type DriverIdKHR = DriverId

pub type ConformanceVersionKHR = ConformanceVersion

pub type PhysicalDeviceDriverPropertiesKHR = PhysicalDeviceDriverProperties



// VK_KHR_shader_float_controls is a preprocessor guard. Do not pass it to API calls.
const khr_shader_float_controls = 1
pub const khr_shader_float_controls_spec_version = 4
pub const khr_shader_float_controls_extension_name = "VK_KHR_shader_float_controls"
pub type ShaderFloatControlsIndependenceKHR = ShaderFloatControlsIndependence

pub type PhysicalDeviceFloatControlsPropertiesKHR = PhysicalDeviceFloatControlsProperties



// VK_KHR_depth_stencil_resolve is a preprocessor guard. Do not pass it to API calls.
const khr_depth_stencil_resolve = 1
pub const khr_depth_stencil_resolve_spec_version = 1
pub const khr_depth_stencil_resolve_extension_name = "VK_KHR_depth_stencil_resolve"
pub type ResolveModeFlagBitsKHR = ResolveModeFlagBits

pub type SubpassDescriptionDepthStencilResolveKHR = SubpassDescriptionDepthStencilResolve

pub type PhysicalDeviceDepthStencilResolvePropertiesKHR = PhysicalDeviceDepthStencilResolveProperties



// VK_KHR_swapchain_mutable_format is a preprocessor guard. Do not pass it to API calls.
const khr_swapchain_mutable_format = 1
pub const khr_swapchain_mutable_format_spec_version = 1
pub const khr_swapchain_mutable_format_extension_name = "VK_KHR_swapchain_mutable_format"


// VK_KHR_timeline_semaphore is a preprocessor guard. Do not pass it to API calls.
const khr_timeline_semaphore = 1
pub const khr_timeline_semaphore_spec_version = 2
pub const khr_timeline_semaphore_extension_name = "VK_KHR_timeline_semaphore"
pub type SemaphoreTypeKHR = SemaphoreType

pub type SemaphoreWaitFlagBitsKHR = SemaphoreWaitFlagBits

pub type PhysicalDeviceTimelineSemaphoreFeaturesKHR = PhysicalDeviceTimelineSemaphoreFeatures

pub type PhysicalDeviceTimelineSemaphorePropertiesKHR = PhysicalDeviceTimelineSemaphoreProperties

pub type SemaphoreTypeCreateInfoKHR = SemaphoreTypeCreateInfo

pub type TimelineSemaphoreSubmitInfoKHR = TimelineSemaphoreSubmitInfo

pub type SemaphoreWaitInfoKHR = SemaphoreWaitInfo

pub type SemaphoreSignalInfoKHR = SemaphoreSignalInfo

type VkGetSemaphoreCounterValueKHR = fn (     C.Device,     C.Semaphore,     &u64) Result

pub fn get_semaphore_counter_value_khr(
    device                                          C.Device,
    semaphore                                       C.Semaphore,
    p_value                                         &u64) Result {
      f := VkGetSemaphoreCounterValueKHR((*loader_p).get_sym('vkGetSemaphoreCounterValueKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetSemaphoreCounterValueKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    semaphore,
    p_value)
}


type VkWaitSemaphoresKHR = fn (     C.Device,     &SemaphoreWaitInfo,     u64) Result

pub fn wait_semaphores_khr(
    device                                          C.Device,
    p_wait_info                                     &SemaphoreWaitInfo,
    timeout                                         u64) Result {
      f := VkWaitSemaphoresKHR((*loader_p).get_sym('vkWaitSemaphoresKHR'
    ) or { 
        println("Couldn't load symbol for 'vkWaitSemaphoresKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_wait_info,
    timeout)
}


type VkSignalSemaphoreKHR = fn (     C.Device,     &SemaphoreSignalInfo) Result

pub fn signal_semaphore_khr(
    device                                          C.Device,
    p_signal_info                                   &SemaphoreSignalInfo) Result {
      f := VkSignalSemaphoreKHR((*loader_p).get_sym('vkSignalSemaphoreKHR'
    ) or { 
        println("Couldn't load symbol for 'vkSignalSemaphoreKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_signal_info)
}




// VK_KHR_vulkan_memory_model is a preprocessor guard. Do not pass it to API calls.
const khr_vulkan_memory_model = 1
pub const khr_vulkan_memory_model_spec_version = 3
pub const khr_vulkan_memory_model_extension_name = "VK_KHR_vulkan_memory_model"
pub type PhysicalDeviceVulkanMemoryModelFeaturesKHR = PhysicalDeviceVulkanMemoryModelFeatures



// VK_KHR_shader_terminate_invocation is a preprocessor guard. Do not pass it to API calls.
const khr_shader_terminate_invocation = 1
pub const khr_shader_terminate_invocation_spec_version = 1
pub const khr_shader_terminate_invocation_extension_name = "VK_KHR_shader_terminate_invocation"
pub type PhysicalDeviceShaderTerminateInvocationFeaturesKHR = PhysicalDeviceShaderTerminateInvocationFeatures



// VK_KHR_fragment_shading_rate is a preprocessor guard. Do not pass it to API calls.
const khr_fragment_shading_rate = 1
pub const khr_fragment_shading_rate_spec_version = 2
pub const khr_fragment_shading_rate_extension_name = "VK_KHR_fragment_shading_rate"

pub enum FragmentShadingRateCombinerOpKHR {
    fragment_shading_rate_combiner_op_keep_khr = int(0)
    fragment_shading_rate_combiner_op_replace_khr = int(1)
    fragment_shading_rate_combiner_op_min_khr = int(2)
    fragment_shading_rate_combiner_op_max_khr = int(3)
    fragment_shading_rate_combiner_op_mul_khr = int(4)
    fragment_shading_rate_combiner_op_max_enum_khr = int(0x7FFFFFFF)
}

// FragmentShadingRateAttachmentInfoKHR extends VkSubpassDescription2
pub struct FragmentShadingRateAttachmentInfoKHR {
mut:
    s_type                               StructureType
    p_next                               voidptr
    p_fragment_shading_rate_attachment   &AttachmentReference2
    shading_rate_attachment_texel_size   Extent2D
} 

// PipelineFragmentShadingRateStateCreateInfoKHR extends VkGraphicsPipelineCreateInfo
pub struct PipelineFragmentShadingRateStateCreateInfoKHR {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    fragment_size                             Extent2D
    combiner_ops                              []FragmentShadingRateCombinerOpKHR
} 

// PhysicalDeviceFragmentShadingRateFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceFragmentShadingRateFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pipeline_fragment_shading_rate Bool32
    primitive_fragment_shading_rate Bool32
    attachment_fragment_shading_rate Bool32
} 

// PhysicalDeviceFragmentShadingRatePropertiesKHR extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceFragmentShadingRatePropertiesKHR {
mut:
    s_type                       StructureType
    p_next                       voidptr
    min_fragment_shading_rate_attachment_texel_size Extent2D
    max_fragment_shading_rate_attachment_texel_size Extent2D
    max_fragment_shading_rate_attachment_texel_size_aspect_ratio u32
    primitive_fragment_shading_rate_with_multiple_viewports Bool32
    layered_shading_rate_attachments Bool32
    fragment_shading_rate_non_trivial_combiner_ops Bool32
    max_fragment_size            Extent2D
    max_fragment_size_aspect_ratio u32
    max_fragment_shading_rate_coverage_samples u32
    max_fragment_shading_rate_rasterization_samples SampleCountFlagBits
    fragment_shading_rate_with_shader_depth_stencil_writes Bool32
    fragment_shading_rate_with_sample_mask Bool32
    fragment_shading_rate_with_shader_sample_mask Bool32
    fragment_shading_rate_with_conservative_rasterization Bool32
    fragment_shading_rate_with_fragment_shader_interlock Bool32
    fragment_shading_rate_with_custom_sample_locations Bool32
    fragment_shading_rate_strict_multiply_combiner Bool32
} 

pub struct PhysicalDeviceFragmentShadingRateKHR {
mut:
    s_type                    StructureType
    p_next                    voidptr
    sample_counts             SampleCountFlags
    fragment_size             Extent2D
} 

type VkGetPhysicalDeviceFragmentShadingRatesKHR = fn (     C.PhysicalDevice,     &u32,     &PhysicalDeviceFragmentShadingRateKHR) Result

pub fn get_physical_device_fragment_shading_rates_khr(
    physical_device                                 C.PhysicalDevice,
    p_fragment_shading_rate_count                   &u32,
    p_fragment_shading_rates                        &PhysicalDeviceFragmentShadingRateKHR) Result {
      f := VkGetPhysicalDeviceFragmentShadingRatesKHR((*loader_p).get_sym('vkGetPhysicalDeviceFragmentShadingRatesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceFragmentShadingRatesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_fragment_shading_rate_count,
    p_fragment_shading_rates)
}


type VkCmdSetFragmentShadingRateKHR = fn (     C.CommandBuffer,     &Extent2D,     []FragmentShadingRateCombinerOpKHR) 

pub fn cmd_set_fragment_shading_rate_khr(
    command_buffer                                  C.CommandBuffer,
    p_fragment_size                                 &Extent2D,
    combiner_ops                                    []FragmentShadingRateCombinerOpKHR)  {
      f := VkCmdSetFragmentShadingRateKHR((*loader_p).get_sym('vkCmdSetFragmentShadingRateKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetFragmentShadingRateKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_fragment_size,
    combiner_ops)
}




// VK_KHR_spirv_1_4 is a preprocessor guard. Do not pass it to API calls.
const khr_spirv_1_4 = 1
pub const khr_spirv_1_4_spec_version        = 1
pub const khr_spirv_1_4_extension_name      = "VK_KHR_spirv_1_4"


// VK_KHR_surface_protected_capabilities is a preprocessor guard. Do not pass it to API calls.
const khr_surface_protected_capabilities = 1
pub const khr_surface_protected_capabilities_spec_version = 1
pub const khr_surface_protected_capabilities_extension_name = "VK_KHR_surface_protected_capabilities"
// SurfaceProtectedCapabilitiesKHR extends VkSurfaceCapabilities2KHR
pub struct SurfaceProtectedCapabilitiesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    supports_protected     Bool32
} 



// VK_KHR_separate_depth_stencil_layouts is a preprocessor guard. Do not pass it to API calls.
const khr_separate_depth_stencil_layouts = 1
pub const khr_separate_depth_stencil_layouts_spec_version = 1
pub const khr_separate_depth_stencil_layouts_extension_name = "VK_KHR_separate_depth_stencil_layouts"
pub type PhysicalDeviceSeparateDepthStencilLayoutsFeaturesKHR = PhysicalDeviceSeparateDepthStencilLayoutsFeatures

pub type AttachmentReferenceStencilLayoutKHR = AttachmentReferenceStencilLayout

pub type AttachmentDescriptionStencilLayoutKHR = AttachmentDescriptionStencilLayout



// VK_KHR_present_wait is a preprocessor guard. Do not pass it to API calls.
const khr_present_wait = 1
pub const khr_present_wait_spec_version     = 1
pub const khr_present_wait_extension_name   = "VK_KHR_present_wait"
// PhysicalDevicePresentWaitFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePresentWaitFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    present_wait           Bool32
} 

type VkWaitForPresentKHR = fn (     C.Device,     C.SwapchainKHR,     u64,     u64) Result

pub fn wait_for_present_khr(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR,
    present_id                                      u64,
    timeout                                         u64) Result {
      f := VkWaitForPresentKHR((*loader_p).get_sym('vkWaitForPresentKHR'
    ) or { 
        println("Couldn't load symbol for 'vkWaitForPresentKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain,
    present_id,
    timeout)
}




// VK_KHR_uniform_buffer_standard_layout is a preprocessor guard. Do not pass it to API calls.
const khr_uniform_buffer_standard_layout = 1
pub const khr_uniform_buffer_standard_layout_spec_version = 1
pub const khr_uniform_buffer_standard_layout_extension_name = "VK_KHR_uniform_buffer_standard_layout"
pub type PhysicalDeviceUniformBufferStandardLayoutFeaturesKHR = PhysicalDeviceUniformBufferStandardLayoutFeatures



// VK_KHR_buffer_device_address is a preprocessor guard. Do not pass it to API calls.
const khr_buffer_device_address = 1
pub const khr_buffer_device_address_spec_version = 1
pub const khr_buffer_device_address_extension_name = "VK_KHR_buffer_device_address"
pub type PhysicalDeviceBufferDeviceAddressFeaturesKHR = PhysicalDeviceBufferDeviceAddressFeatures

pub type BufferDeviceAddressInfoKHR = BufferDeviceAddressInfo

pub type BufferOpaqueCaptureAddressCreateInfoKHR = BufferOpaqueCaptureAddressCreateInfo

pub type MemoryOpaqueCaptureAddressAllocateInfoKHR = MemoryOpaqueCaptureAddressAllocateInfo

pub type DeviceMemoryOpaqueCaptureAddressInfoKHR = DeviceMemoryOpaqueCaptureAddressInfo

type VkGetBufferDeviceAddressKHR = fn (     C.Device,     &BufferDeviceAddressInfo) DeviceAddress

pub fn get_buffer_device_address_khr(
    device                                          C.Device,
    p_info                                          &BufferDeviceAddressInfo) DeviceAddress {
      f := VkGetBufferDeviceAddressKHR((*loader_p).get_sym("vkGetBufferDeviceAddressKHR"
    ) or { 
        panic("Couldn't load symbol for 'vkGetBufferDeviceAddressKHR': ${err}") })
    return f(
    device,
    p_info)
}


type VkGetBufferOpaqueCaptureAddressKHR = fn (     C.Device,     &BufferDeviceAddressInfo) u64

pub fn get_buffer_opaque_capture_address_khr(
    device                                          C.Device,
    p_info                                          &BufferDeviceAddressInfo) u64 {
      f := VkGetBufferOpaqueCaptureAddressKHR((*loader_p).get_sym("vkGetBufferOpaqueCaptureAddressKHR"
    ) or { 
        panic("Couldn't load symbol for 'vkGetBufferOpaqueCaptureAddressKHR': ${err}") })
    return f(
    device,
    p_info)
}


type VkGetDeviceMemoryOpaqueCaptureAddressKHR = fn (     C.Device,     &DeviceMemoryOpaqueCaptureAddressInfo) u64

pub fn get_device_memory_opaque_capture_address_khr(
    device                                          C.Device,
    p_info                                          &DeviceMemoryOpaqueCaptureAddressInfo) u64 {
      f := VkGetDeviceMemoryOpaqueCaptureAddressKHR((*loader_p).get_sym("vkGetDeviceMemoryOpaqueCaptureAddressKHR"
    ) or { 
        panic("Couldn't load symbol for 'vkGetDeviceMemoryOpaqueCaptureAddressKHR': ${err}") })
    return f(
    device,
    p_info)
}




// VK_KHR_deferred_host_operations is a preprocessor guard. Do not pass it to API calls.
const khr_deferred_host_operations = 1
pub type C.DeferredOperationKHR = voidptr
pub const khr_deferred_host_operations_spec_version = 4
pub const khr_deferred_host_operations_extension_name = "VK_KHR_deferred_host_operations"
type VkCreateDeferredOperationKHR = fn (     C.Device,     &AllocationCallbacks,     &C.DeferredOperationKHR) Result

pub fn create_deferred_operation_khr(
    device                                          C.Device,
    p_allocator                                     &AllocationCallbacks,
    p_deferred_operation                            &C.DeferredOperationKHR) Result {
      f := VkCreateDeferredOperationKHR((*loader_p).get_sym('vkCreateDeferredOperationKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateDeferredOperationKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_allocator,
    p_deferred_operation)
}


type VkDestroyDeferredOperationKHR = fn (     C.Device,     C.DeferredOperationKHR,     &AllocationCallbacks) 

pub fn destroy_deferred_operation_khr(
    device                                          C.Device,
    operation                                       C.DeferredOperationKHR,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyDeferredOperationKHR((*loader_p).get_sym('vkDestroyDeferredOperationKHR'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyDeferredOperationKHR': ${err}")
        return 
    })
    f(
    device,
    operation,
    p_allocator)
}


type VkGetDeferredOperationMaxConcurrencyKHR = fn (     C.Device,     C.DeferredOperationKHR) u32

pub fn get_deferred_operation_max_concurrency_khr(
    device                                          C.Device,
    operation                                       C.DeferredOperationKHR) u32 {
      f := VkGetDeferredOperationMaxConcurrencyKHR((*loader_p).get_sym("vkGetDeferredOperationMaxConcurrencyKHR"
    ) or { 
        panic("Couldn't load symbol for 'vkGetDeferredOperationMaxConcurrencyKHR': ${err}") })
    return f(
    device,
    operation)
}


type VkGetDeferredOperationResultKHR = fn (     C.Device,     C.DeferredOperationKHR) Result

pub fn get_deferred_operation_result_khr(
    device                                          C.Device,
    operation                                       C.DeferredOperationKHR) Result {
      f := VkGetDeferredOperationResultKHR((*loader_p).get_sym('vkGetDeferredOperationResultKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeferredOperationResultKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    operation)
}


type VkDeferredOperationJoinKHR = fn (     C.Device,     C.DeferredOperationKHR) Result

pub fn deferred_operation_join_khr(
    device                                          C.Device,
    operation                                       C.DeferredOperationKHR) Result {
      f := VkDeferredOperationJoinKHR((*loader_p).get_sym('vkDeferredOperationJoinKHR'
    ) or { 
        println("Couldn't load symbol for 'vkDeferredOperationJoinKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    operation)
}




// VK_KHR_pipeline_executable_properties is a preprocessor guard. Do not pass it to API calls.
const khr_pipeline_executable_properties = 1
pub const khr_pipeline_executable_properties_spec_version = 1
pub const khr_pipeline_executable_properties_extension_name = "VK_KHR_pipeline_executable_properties"

pub enum PipelineExecutableStatisticFormatKHR {
    pipeline_executable_statistic_format_bool32_khr = int(0)
    pipeline_executable_statistic_format_int64_khr = int(1)
    pipeline_executable_statistic_format_uint64_khr = int(2)
    pipeline_executable_statistic_format_float64_khr = int(3)
    pipeline_executable_statistic_format_max_enum_khr = int(0x7FFFFFFF)
}

// PhysicalDevicePipelineExecutablePropertiesFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePipelineExecutablePropertiesFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pipeline_executable_info Bool32
} 

pub struct PipelineInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pipeline               C.Pipeline
} 

pub struct PipelineExecutablePropertiesKHR {
mut:
    s_type                    StructureType
    p_next                    voidptr
    stages                    ShaderStageFlags
    name                      []char
    description               []char
    subgroup_size             u32
} 

pub struct PipelineExecutableInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pipeline               C.Pipeline
    executable_index       u32
} 

pub union PipelineExecutableStatisticValueKHR {
mut:
    b32             Bool32
    i64             i64
    u64             u64
    f64             f64
} 

pub struct PipelineExecutableStatisticKHR {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    name                                          []char
    description                                   []char
    format                                        PipelineExecutableStatisticFormatKHR
    value                                         PipelineExecutableStatisticValueKHR
} 

pub struct PipelineExecutableInternalRepresentationKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    name                   []char
    description            []char
    is_text                Bool32
    data_size              usize
    p_data                 voidptr
} 

type VkGetPipelineExecutablePropertiesKHR = fn (     C.Device,     &PipelineInfoKHR,     &u32,     &PipelineExecutablePropertiesKHR) Result

pub fn get_pipeline_executable_properties_khr(
    device                                          C.Device,
    p_pipeline_info                                 &PipelineInfoKHR,
    p_executable_count                              &u32,
    p_properties                                    &PipelineExecutablePropertiesKHR) Result {
      f := VkGetPipelineExecutablePropertiesKHR((*loader_p).get_sym('vkGetPipelineExecutablePropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPipelineExecutablePropertiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_pipeline_info,
    p_executable_count,
    p_properties)
}


type VkGetPipelineExecutableStatisticsKHR = fn (     C.Device,     &PipelineExecutableInfoKHR,     &u32,     &PipelineExecutableStatisticKHR) Result

pub fn get_pipeline_executable_statistics_khr(
    device                                          C.Device,
    p_executable_info                               &PipelineExecutableInfoKHR,
    p_statistic_count                               &u32,
    p_statistics                                    &PipelineExecutableStatisticKHR) Result {
      f := VkGetPipelineExecutableStatisticsKHR((*loader_p).get_sym('vkGetPipelineExecutableStatisticsKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPipelineExecutableStatisticsKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_executable_info,
    p_statistic_count,
    p_statistics)
}


type VkGetPipelineExecutableInternalRepresentationsKHR = fn (     C.Device,     &PipelineExecutableInfoKHR,     &u32,     &PipelineExecutableInternalRepresentationKHR) Result

pub fn get_pipeline_executable_internal_representations_khr(
    device                                          C.Device,
    p_executable_info                               &PipelineExecutableInfoKHR,
    p_internal_representation_count                 &u32,
    p_internal_representations                      &PipelineExecutableInternalRepresentationKHR) Result {
      f := VkGetPipelineExecutableInternalRepresentationsKHR((*loader_p).get_sym('vkGetPipelineExecutableInternalRepresentationsKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPipelineExecutableInternalRepresentationsKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_executable_info,
    p_internal_representation_count,
    p_internal_representations)
}




// VK_KHR_map_memory2 is a preprocessor guard. Do not pass it to API calls.
const khr_map_memory2 = 1
pub const khr_map_memory_2_spec_version     = 1
pub const khr_map_memory_2_extension_name   = "VK_KHR_map_memory2"
pub type MemoryUnmapFlagsKHR = u32
pub struct MemoryMapInfoKHR {
mut:
    s_type                  StructureType
    p_next                  voidptr
    flags                   MemoryMapFlags
    memory                  C.DeviceMemory
    offset                  DeviceSize
    size                    DeviceSize
} 

pub struct MemoryUnmapInfoKHR {
mut:
    s_type                       StructureType
    p_next                       voidptr
    flags                        MemoryUnmapFlagsKHR
    memory                       C.DeviceMemory
} 

type VkMapMemory2KHR = fn (     C.Device,     &MemoryMapInfoKHR,     &voidptr) Result

pub fn map_memory2_khr(
    device                                          C.Device,
    p_memory_map_info                               &MemoryMapInfoKHR,
    pp_data                                         &voidptr) Result {
      f := VkMapMemory2KHR((*loader_p).get_sym('vkMapMemory2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkMapMemory2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_memory_map_info,
    pp_data)
}


type VkUnmapMemory2KHR = fn (     C.Device,     &MemoryUnmapInfoKHR) Result

pub fn unmap_memory2_khr(
    device                                          C.Device,
    p_memory_unmap_info                             &MemoryUnmapInfoKHR) Result {
      f := VkUnmapMemory2KHR((*loader_p).get_sym('vkUnmapMemory2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkUnmapMemory2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_memory_unmap_info)
}




// VK_KHR_shader_integer_dot_product is a preprocessor guard. Do not pass it to API calls.
const khr_shader_integer_dot_product = 1
pub const khr_shader_integer_dot_product_spec_version = 1
pub const khr_shader_integer_dot_product_extension_name = "VK_KHR_shader_integer_dot_product"
pub type PhysicalDeviceShaderIntegerDotProductFeaturesKHR = PhysicalDeviceShaderIntegerDotProductFeatures

pub type PhysicalDeviceShaderIntegerDotProductPropertiesKHR = PhysicalDeviceShaderIntegerDotProductProperties



// VK_KHR_pipeline_library is a preprocessor guard. Do not pass it to API calls.
const khr_pipeline_library = 1
pub const khr_pipeline_library_spec_version = 1
pub const khr_pipeline_library_extension_name = "VK_KHR_pipeline_library"
// PipelineLibraryCreateInfoKHR extends VkGraphicsPipelineCreateInfo
pub struct PipelineLibraryCreateInfoKHR {
mut:
    s_type                   StructureType
    p_next                   voidptr
    library_count            u32
    p_libraries              &C.Pipeline
} 



// VK_KHR_shader_non_semantic_info is a preprocessor guard. Do not pass it to API calls.
const khr_shader_non_semantic_info = 1
pub const khr_shader_non_semantic_info_spec_version = 1
pub const khr_shader_non_semantic_info_extension_name = "VK_KHR_shader_non_semantic_info"


// VK_KHR_present_id is a preprocessor guard. Do not pass it to API calls.
const khr_present_id = 1
pub const khr_present_id_spec_version       = 1
pub const khr_present_id_extension_name     = "VK_KHR_present_id"
// PresentIdKHR extends VkPresentInfoKHR
pub struct PresentIdKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    swapchain_count        u32
    p_present_ids          &u64
} 

// PhysicalDevicePresentIdFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePresentIdFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    present_id             Bool32
} 



// VK_KHR_video_encode_queue is a preprocessor guard. Do not pass it to API calls.
const khr_video_encode_queue = 1
pub const khr_video_encode_queue_spec_version = 10
pub const khr_video_encode_queue_extension_name = "VK_KHR_video_encode_queue"

pub enum VideoEncodeTuningModeKHR {
    video_encode_tuning_mode_default_khr = int(0)
    video_encode_tuning_mode_high_quality_khr = int(1)
    video_encode_tuning_mode_low_latency_khr = int(2)
    video_encode_tuning_mode_ultra_low_latency_khr = int(3)
    video_encode_tuning_mode_lossless_khr = int(4)
    video_encode_tuning_mode_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoEncodeFlagsKHR = u32

pub enum VideoEncodeCapabilityFlagBitsKHR {
    video_encode_capability_preceding_externally_encoded_bytes_bit_khr = int(0x00000001)
    video_encode_capability_insufficient_bitstream_buffer_range_detection_bit_khr = int(0x00000002)
    video_encode_capability_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoEncodeCapabilityFlagsKHR = u32

pub enum VideoEncodeRateControlModeFlagBitsKHR {
    video_encode_rate_control_mode_default_khr = int(0)
    video_encode_rate_control_mode_disabled_bit_khr = int(0x00000001)
    video_encode_rate_control_mode_cbr_bit_khr = int(0x00000002)
    video_encode_rate_control_mode_vbr_bit_khr = int(0x00000004)
    video_encode_rate_control_mode_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoEncodeRateControlModeFlagsKHR = u32

pub enum VideoEncodeFeedbackFlagBitsKHR {
    video_encode_feedback_bitstream_buffer_offset_bit_khr = int(0x00000001)
    video_encode_feedback_bitstream_bytes_written_bit_khr = int(0x00000002)
    video_encode_feedback_bitstream_has_overrides_bit_khr = int(0x00000004)
    video_encode_feedback_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoEncodeFeedbackFlagsKHR = u32

pub enum VideoEncodeUsageFlagBitsKHR {
    video_encode_usage_default_khr = int(0)
    video_encode_usage_transcoding_bit_khr = int(0x00000001)
    video_encode_usage_streaming_bit_khr = int(0x00000002)
    video_encode_usage_recording_bit_khr = int(0x00000004)
    video_encode_usage_conferencing_bit_khr = int(0x00000008)
    video_encode_usage_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoEncodeUsageFlagsKHR = u32

pub enum VideoEncodeContentFlagBitsKHR {
    video_encode_content_default_khr = int(0)
    video_encode_content_camera_bit_khr = int(0x00000001)
    video_encode_content_desktop_bit_khr = int(0x00000002)
    video_encode_content_rendered_bit_khr = int(0x00000004)
    video_encode_content_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type VideoEncodeContentFlagsKHR = u32
pub type VideoEncodeRateControlFlagsKHR = u32
pub struct VideoEncodeInfoKHR {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    flags                                     VideoEncodeFlagsKHR
    dst_buffer                                C.Buffer
    dst_buffer_offset                         DeviceSize
    dst_buffer_range                          DeviceSize
    src_picture_resource                      VideoPictureResourceInfoKHR
    p_setup_reference_slot                    &VideoReferenceSlotInfoKHR
    reference_slot_count                      u32
    p_reference_slots                         &VideoReferenceSlotInfoKHR
    preceding_externally_encoded_bytes        u32
} 

// VideoEncodeCapabilitiesKHR extends VkVideoCapabilitiesKHR
pub struct VideoEncodeCapabilitiesKHR {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    flags                                       VideoEncodeCapabilityFlagsKHR
    rate_control_modes                          VideoEncodeRateControlModeFlagsKHR
    max_rate_control_layers                     u32
    max_bitrate                                 u64
    max_quality_levels                          u32
    encode_input_picture_granularity            Extent2D
    supported_encode_feedback_flags             VideoEncodeFeedbackFlagsKHR
} 

// QueryPoolVideoEncodeFeedbackCreateInfoKHR extends VkQueryPoolCreateInfo
pub struct QueryPoolVideoEncodeFeedbackCreateInfoKHR {
mut:
    s_type                               StructureType
    p_next                               voidptr
    encode_feedback_flags                VideoEncodeFeedbackFlagsKHR
} 

// VideoEncodeUsageInfoKHR extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub struct VideoEncodeUsageInfoKHR {
mut:
    s_type                              StructureType
    p_next                              voidptr
    video_usage_hints                   VideoEncodeUsageFlagsKHR
    video_content_hints                 VideoEncodeContentFlagsKHR
    tuning_mode                         VideoEncodeTuningModeKHR
} 

pub struct VideoEncodeRateControlLayerInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    average_bitrate        u64
    max_bitrate            u64
    frame_rate_numerator   u32
    frame_rate_denominator u32
} 

// VideoEncodeRateControlInfoKHR extends VkVideoCodingControlInfoKHR,VkVideoBeginCodingInfoKHR
pub struct VideoEncodeRateControlInfoKHR {
mut:
    s_type                                             StructureType
    p_next                                             voidptr
    flags                                              VideoEncodeRateControlFlagsKHR
    rate_control_mode                                  VideoEncodeRateControlModeFlagBitsKHR
    layer_count                                        u32
    p_layers                                           &VideoEncodeRateControlLayerInfoKHR
    virtual_buffer_size_in_ms                          u32
    initial_virtual_buffer_size_in_ms                  u32
} 

pub struct PhysicalDeviceVideoEncodeQualityLevelInfoKHR {
mut:
    s_type                              StructureType
    p_next                              voidptr
    p_video_profile                     &VideoProfileInfoKHR
    quality_level                       u32
} 

pub struct VideoEncodeQualityLevelPropertiesKHR {
mut:
    s_type                                         StructureType
    p_next                                         voidptr
    preferred_rate_control_mode                    VideoEncodeRateControlModeFlagBitsKHR
    preferred_rate_control_layer_count             u32
} 

// VideoEncodeQualityLevelInfoKHR extends VkVideoCodingControlInfoKHR,VkVideoSessionParametersCreateInfoKHR
pub struct VideoEncodeQualityLevelInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    quality_level          u32
} 

pub struct VideoEncodeSessionParametersGetInfoKHR {
mut:
    s_type                             StructureType
    p_next                             voidptr
    video_session_parameters           C.VideoSessionParametersKHR
} 

pub struct VideoEncodeSessionParametersFeedbackInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    has_overrides          Bool32
} 

type VkGetPhysicalDeviceVideoEncodeQualityLevelPropertiesKHR = fn (     C.PhysicalDevice,     &PhysicalDeviceVideoEncodeQualityLevelInfoKHR,     &VideoEncodeQualityLevelPropertiesKHR) Result

pub fn get_physical_device_video_encode_quality_level_properties_khr(
    physical_device                                 C.PhysicalDevice,
    p_quality_level_info                            &PhysicalDeviceVideoEncodeQualityLevelInfoKHR,
    p_quality_level_properties                      &VideoEncodeQualityLevelPropertiesKHR) Result {
      f := VkGetPhysicalDeviceVideoEncodeQualityLevelPropertiesKHR((*loader_p).get_sym('vkGetPhysicalDeviceVideoEncodeQualityLevelPropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceVideoEncodeQualityLevelPropertiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_quality_level_info,
    p_quality_level_properties)
}


type VkGetEncodedVideoSessionParametersKHR = fn (     C.Device,     &VideoEncodeSessionParametersGetInfoKHR,     &VideoEncodeSessionParametersFeedbackInfoKHR,     &usize,     voidptr) Result

pub fn get_encoded_video_session_parameters_khr(
    device                                          C.Device,
    p_video_session_parameters_info                 &VideoEncodeSessionParametersGetInfoKHR,
    p_feedback_info                                 &VideoEncodeSessionParametersFeedbackInfoKHR,
    p_data_size                                     &usize,
    p_data                                          voidptr) Result {
      f := VkGetEncodedVideoSessionParametersKHR((*loader_p).get_sym('vkGetEncodedVideoSessionParametersKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetEncodedVideoSessionParametersKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_video_session_parameters_info,
    p_feedback_info,
    p_data_size,
    p_data)
}


type VkCmdEncodeVideoKHR = fn (     C.CommandBuffer,     &VideoEncodeInfoKHR) 

pub fn cmd_encode_video_khr(
    command_buffer                                  C.CommandBuffer,
    p_encode_info                                   &VideoEncodeInfoKHR)  {
      f := VkCmdEncodeVideoKHR((*loader_p).get_sym('vkCmdEncodeVideoKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEncodeVideoKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_encode_info)
}




// VK_KHR_synchronization2 is a preprocessor guard. Do not pass it to API calls.
const khr_synchronization2 = 1
pub const khr_synchronization_2_spec_version = 1
pub const khr_synchronization_2_extension_name = "VK_KHR_synchronization2"
pub type PipelineStageFlagBits2KHR = u64

pub type AccessFlagBits2KHR = u64

pub type SubmitFlagBitsKHR = SubmitFlagBits

pub type MemoryBarrier2KHR = MemoryBarrier2

pub type BufferMemoryBarrier2KHR = BufferMemoryBarrier2

pub type ImageMemoryBarrier2KHR = ImageMemoryBarrier2

pub type DependencyInfoKHR = DependencyInfo

pub type SubmitInfo2KHR = SubmitInfo2

pub type SemaphoreSubmitInfoKHR = SemaphoreSubmitInfo

pub type CommandBufferSubmitInfoKHR = CommandBufferSubmitInfo

pub type PhysicalDeviceSynchronization2FeaturesKHR = PhysicalDeviceSynchronization2Features

// QueueFamilyCheckpointProperties2NV extends VkQueueFamilyProperties2
pub struct QueueFamilyCheckpointProperties2NV {
mut:
    s_type                       StructureType
    p_next                       voidptr
    checkpoint_execution_stage_mask PipelineStageFlags2
} 

pub struct CheckpointData2NV {
mut:
    s_type                       StructureType
    p_next                       voidptr
    stage                        PipelineStageFlags2
    p_checkpoint_marker          voidptr
} 

type VkCmdSetEvent2KHR = fn (     C.CommandBuffer,     C.Event,     &DependencyInfo) 

pub fn cmd_set_event2_khr(
    command_buffer                                  C.CommandBuffer,
    event                                           C.Event,
    p_dependency_info                               &DependencyInfo)  {
      f := VkCmdSetEvent2KHR((*loader_p).get_sym('vkCmdSetEvent2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetEvent2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    event,
    p_dependency_info)
}


type VkCmdResetEvent2KHR = fn (     C.CommandBuffer,     C.Event,     PipelineStageFlags2) 

pub fn cmd_reset_event2_khr(
    command_buffer                                  C.CommandBuffer,
    event                                           C.Event,
    stage_mask                                      PipelineStageFlags2)  {
      f := VkCmdResetEvent2KHR((*loader_p).get_sym('vkCmdResetEvent2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdResetEvent2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    event,
    stage_mask)
}


type VkCmdWaitEvents2KHR = fn (     C.CommandBuffer,     u32,     &C.Event,     &DependencyInfo) 

pub fn cmd_wait_events2_khr(
    command_buffer                                  C.CommandBuffer,
    event_count                                     u32,
    p_events                                        &C.Event,
    p_dependency_infos                              &DependencyInfo)  {
      f := VkCmdWaitEvents2KHR((*loader_p).get_sym('vkCmdWaitEvents2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdWaitEvents2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    event_count,
    p_events,
    p_dependency_infos)
}


type VkCmdPipelineBarrier2KHR = fn (     C.CommandBuffer,     &DependencyInfo) 

pub fn cmd_pipeline_barrier2_khr(
    command_buffer                                  C.CommandBuffer,
    p_dependency_info                               &DependencyInfo)  {
      f := VkCmdPipelineBarrier2KHR((*loader_p).get_sym('vkCmdPipelineBarrier2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdPipelineBarrier2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_dependency_info)
}


type VkCmdWriteTimestamp2KHR = fn (     C.CommandBuffer,     PipelineStageFlags2,     C.QueryPool,     u32) 

pub fn cmd_write_timestamp2_khr(
    command_buffer                                  C.CommandBuffer,
    stage                                           PipelineStageFlags2,
    query_pool                                      C.QueryPool,
    query                                           u32)  {
      f := VkCmdWriteTimestamp2KHR((*loader_p).get_sym('vkCmdWriteTimestamp2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdWriteTimestamp2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    stage,
    query_pool,
    query)
}


type VkQueueSubmit2KHR = fn (     C.Queue,     u32,     &SubmitInfo2,     C.Fence) Result

pub fn queue_submit2_khr(
    queue                                           C.Queue,
    submit_count                                    u32,
    p_submits                                       &SubmitInfo2,
    fence                                           C.Fence) Result {
      f := VkQueueSubmit2KHR((*loader_p).get_sym('vkQueueSubmit2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkQueueSubmit2KHR': ${err}")
        return Result.error_unknown
    })
    return f(
    queue,
    submit_count,
    p_submits,
    fence)
}


type VkCmdWriteBufferMarker2AMD = fn (     C.CommandBuffer,     PipelineStageFlags2,     C.Buffer,     DeviceSize,     u32) 

pub fn cmd_write_buffer_marker2_amd(
    command_buffer                                  C.CommandBuffer,
    stage                                           PipelineStageFlags2,
    dst_buffer                                      C.Buffer,
    dst_offset                                      DeviceSize,
    marker                                          u32)  {
      f := VkCmdWriteBufferMarker2AMD((*loader_p).get_sym('vkCmdWriteBufferMarker2AMD'
    ) or { 
        println("Couldn't load symbol for 'vkCmdWriteBufferMarker2AMD': ${err}")
        return 
    })
    f(
    command_buffer,
    stage,
    dst_buffer,
    dst_offset,
    marker)
}


type VkGetQueueCheckpointData2NV = fn (     C.Queue,     &u32,     &CheckpointData2NV) 

pub fn get_queue_checkpoint_data2_nv(
    queue                                           C.Queue,
    p_checkpoint_data_count                         &u32,
    p_checkpoint_data                               &CheckpointData2NV)  {
      f := VkGetQueueCheckpointData2NV((*loader_p).get_sym('vkGetQueueCheckpointData2NV'
    ) or { 
        println("Couldn't load symbol for 'vkGetQueueCheckpointData2NV': ${err}")
        return 
    })
    f(
    queue,
    p_checkpoint_data_count,
    p_checkpoint_data)
}




// VK_KHR_fragment_shader_barycentric is a preprocessor guard. Do not pass it to API calls.
const khr_fragment_shader_barycentric = 1
pub const khr_fragment_shader_barycentric_spec_version = 1
pub const khr_fragment_shader_barycentric_extension_name = "VK_KHR_fragment_shader_barycentric"
// PhysicalDeviceFragmentShaderBarycentricFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceFragmentShaderBarycentricFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    fragment_shader_barycentric Bool32
} 

// PhysicalDeviceFragmentShaderBarycentricPropertiesKHR extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceFragmentShaderBarycentricPropertiesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    tri_strip_vertex_order_independent_of_provoking_vertex Bool32
} 



// VK_KHR_shader_subgroup_uniform_control_flow is a preprocessor guard. Do not pass it to API calls.
const khr_shader_subgroup_uniform_control_flow = 1
pub const khr_shader_subgroup_uniform_control_flow_spec_version = 1
pub const khr_shader_subgroup_uniform_control_flow_extension_name = "VK_KHR_shader_subgroup_uniform_control_flow"
// PhysicalDeviceShaderSubgroupUniformControlFlowFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderSubgroupUniformControlFlowFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_subgroup_uniform_control_flow Bool32
} 



// VK_KHR_zero_initialize_workgroup_memory is a preprocessor guard. Do not pass it to API calls.
const khr_zero_initialize_workgroup_memory = 1
pub const khr_zero_initialize_workgroup_memory_spec_version = 1
pub const khr_zero_initialize_workgroup_memory_extension_name = "VK_KHR_zero_initialize_workgroup_memory"
pub type PhysicalDeviceZeroInitializeWorkgroupMemoryFeaturesKHR = PhysicalDeviceZeroInitializeWorkgroupMemoryFeatures



// VK_KHR_workgroup_memory_explicit_layout is a preprocessor guard. Do not pass it to API calls.
const khr_workgroup_memory_explicit_layout = 1
pub const khr_workgroup_memory_explicit_layout_spec_version = 1
pub const khr_workgroup_memory_explicit_layout_extension_name = "VK_KHR_workgroup_memory_explicit_layout"
// PhysicalDeviceWorkgroupMemoryExplicitLayoutFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceWorkgroupMemoryExplicitLayoutFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    workgroup_memory_explicit_layout Bool32
    workgroup_memory_explicit_layout_scalar_block_layout Bool32
    workgroup_memory_explicit_layout8_bit_access Bool32
    workgroup_memory_explicit_layout16_bit_access Bool32
} 



// VK_KHR_copy_commands2 is a preprocessor guard. Do not pass it to API calls.
const khr_copy_commands2 = 1
pub const khr_copy_commands_2_spec_version  = 1
pub const khr_copy_commands_2_extension_name = "VK_KHR_copy_commands2"
pub type CopyBufferInfo2KHR = CopyBufferInfo2

pub type CopyImageInfo2KHR = CopyImageInfo2

pub type CopyBufferToImageInfo2KHR = CopyBufferToImageInfo2

pub type CopyImageToBufferInfo2KHR = CopyImageToBufferInfo2

pub type BlitImageInfo2KHR = BlitImageInfo2

pub type ResolveImageInfo2KHR = ResolveImageInfo2

pub type BufferCopy2KHR = BufferCopy2

pub type ImageCopy2KHR = ImageCopy2

pub type ImageBlit2KHR = ImageBlit2

pub type BufferImageCopy2KHR = BufferImageCopy2

pub type ImageResolve2KHR = ImageResolve2

type VkCmdCopyBuffer2KHR = fn (     C.CommandBuffer,     &CopyBufferInfo2) 

pub fn cmd_copy_buffer2_khr(
    command_buffer                                  C.CommandBuffer,
    p_copy_buffer_info                              &CopyBufferInfo2)  {
      f := VkCmdCopyBuffer2KHR((*loader_p).get_sym('vkCmdCopyBuffer2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyBuffer2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_copy_buffer_info)
}


type VkCmdCopyImage2KHR = fn (     C.CommandBuffer,     &CopyImageInfo2) 

pub fn cmd_copy_image2_khr(
    command_buffer                                  C.CommandBuffer,
    p_copy_image_info                               &CopyImageInfo2)  {
      f := VkCmdCopyImage2KHR((*loader_p).get_sym('vkCmdCopyImage2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyImage2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_copy_image_info)
}


type VkCmdCopyBufferToImage2KHR = fn (     C.CommandBuffer,     &CopyBufferToImageInfo2) 

pub fn cmd_copy_buffer_to_image2_khr(
    command_buffer                                  C.CommandBuffer,
    p_copy_buffer_to_image_info                     &CopyBufferToImageInfo2)  {
      f := VkCmdCopyBufferToImage2KHR((*loader_p).get_sym('vkCmdCopyBufferToImage2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyBufferToImage2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_copy_buffer_to_image_info)
}


type VkCmdCopyImageToBuffer2KHR = fn (     C.CommandBuffer,     &CopyImageToBufferInfo2) 

pub fn cmd_copy_image_to_buffer2_khr(
    command_buffer                                  C.CommandBuffer,
    p_copy_image_to_buffer_info                     &CopyImageToBufferInfo2)  {
      f := VkCmdCopyImageToBuffer2KHR((*loader_p).get_sym('vkCmdCopyImageToBuffer2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyImageToBuffer2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_copy_image_to_buffer_info)
}


type VkCmdBlitImage2KHR = fn (     C.CommandBuffer,     &BlitImageInfo2) 

pub fn cmd_blit_image2_khr(
    command_buffer                                  C.CommandBuffer,
    p_blit_image_info                               &BlitImageInfo2)  {
      f := VkCmdBlitImage2KHR((*loader_p).get_sym('vkCmdBlitImage2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBlitImage2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_blit_image_info)
}


type VkCmdResolveImage2KHR = fn (     C.CommandBuffer,     &ResolveImageInfo2) 

pub fn cmd_resolve_image2_khr(
    command_buffer                                  C.CommandBuffer,
    p_resolve_image_info                            &ResolveImageInfo2)  {
      f := VkCmdResolveImage2KHR((*loader_p).get_sym('vkCmdResolveImage2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdResolveImage2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_resolve_image_info)
}




// VK_KHR_format_feature_flags2 is a preprocessor guard. Do not pass it to API calls.
const khr_format_feature_flags2 = 1
pub const khr_format_feature_flags_2_spec_version = 2
pub const khr_format_feature_flags_2_extension_name = "VK_KHR_format_feature_flags2"
pub type FormatFeatureFlagBits2KHR = u64

pub type FormatProperties3KHR = FormatProperties3



// VK_KHR_ray_tracing_maintenance1 is a preprocessor guard. Do not pass it to API calls.
const khr_ray_tracing_maintenance1 = 1
pub const khr_ray_tracing_maintenance_1_spec_version = 1
pub const khr_ray_tracing_maintenance_1_extension_name = "VK_KHR_ray_tracing_maintenance1"
// PhysicalDeviceRayTracingMaintenance1FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRayTracingMaintenance1FeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    ray_tracing_maintenance1 Bool32
    ray_tracing_pipeline_trace_rays_indirect2 Bool32
} 

pub struct TraceRaysIndirectCommand2KHR {
mut:
    raygen_shader_record_address DeviceAddress
    raygen_shader_record_size DeviceSize
    miss_shader_binding_table_address DeviceAddress
    miss_shader_binding_table_size DeviceSize
    miss_shader_binding_table_stride DeviceSize
    hit_shader_binding_table_address DeviceAddress
    hit_shader_binding_table_size DeviceSize
    hit_shader_binding_table_stride DeviceSize
    callable_shader_binding_table_address DeviceAddress
    callable_shader_binding_table_size DeviceSize
    callable_shader_binding_table_stride DeviceSize
    width                  u32
    height                 u32
    depth                  u32
} 

type VkCmdTraceRaysIndirect2KHR = fn (     C.CommandBuffer,     DeviceAddress) 

pub fn cmd_trace_rays_indirect2_khr(
    command_buffer                                  C.CommandBuffer,
    indirect_device_address                         DeviceAddress)  {
      f := VkCmdTraceRaysIndirect2KHR((*loader_p).get_sym('vkCmdTraceRaysIndirect2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdTraceRaysIndirect2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    indirect_device_address)
}




// VK_KHR_portability_enumeration is a preprocessor guard. Do not pass it to API calls.
const khr_portability_enumeration = 1
pub const khr_portability_enumeration_spec_version = 1
pub const khr_portability_enumeration_extension_name = "VK_KHR_portability_enumeration"


// VK_KHR_maintenance4 is a preprocessor guard. Do not pass it to API calls.
const khr_maintenance4 = 1
pub const khr_maintenance_4_spec_version    = 2
pub const khr_maintenance_4_extension_name  = "VK_KHR_maintenance4"
pub type PhysicalDeviceMaintenance4FeaturesKHR = PhysicalDeviceMaintenance4Features

pub type PhysicalDeviceMaintenance4PropertiesKHR = PhysicalDeviceMaintenance4Properties

pub type DeviceBufferMemoryRequirementsKHR = DeviceBufferMemoryRequirements

pub type DeviceImageMemoryRequirementsKHR = DeviceImageMemoryRequirements

type VkGetDeviceBufferMemoryRequirementsKHR = fn (     C.Device,     &DeviceBufferMemoryRequirements,     &MemoryRequirements2) 

pub fn get_device_buffer_memory_requirements_khr(
    device                                          C.Device,
    p_info                                          &DeviceBufferMemoryRequirements,
    p_memory_requirements                           &MemoryRequirements2)  {
      f := VkGetDeviceBufferMemoryRequirementsKHR((*loader_p).get_sym('vkGetDeviceBufferMemoryRequirementsKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceBufferMemoryRequirementsKHR': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_memory_requirements)
}


type VkGetDeviceImageMemoryRequirementsKHR = fn (     C.Device,     &DeviceImageMemoryRequirements,     &MemoryRequirements2) 

pub fn get_device_image_memory_requirements_khr(
    device                                          C.Device,
    p_info                                          &DeviceImageMemoryRequirements,
    p_memory_requirements                           &MemoryRequirements2)  {
      f := VkGetDeviceImageMemoryRequirementsKHR((*loader_p).get_sym('vkGetDeviceImageMemoryRequirementsKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceImageMemoryRequirementsKHR': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_memory_requirements)
}


type VkGetDeviceImageSparseMemoryRequirementsKHR = fn (     C.Device,     &DeviceImageMemoryRequirements,     &u32,     &SparseImageMemoryRequirements2) 

pub fn get_device_image_sparse_memory_requirements_khr(
    device                                          C.Device,
    p_info                                          &DeviceImageMemoryRequirements,
    p_sparse_memory_requirement_count               &u32,
    p_sparse_memory_requirements                    &SparseImageMemoryRequirements2)  {
      f := VkGetDeviceImageSparseMemoryRequirementsKHR((*loader_p).get_sym('vkGetDeviceImageSparseMemoryRequirementsKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceImageSparseMemoryRequirementsKHR': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_sparse_memory_requirement_count,
    p_sparse_memory_requirements)
}




// VK_KHR_maintenance5 is a preprocessor guard. Do not pass it to API calls.
const khr_maintenance5 = 1
pub const khr_maintenance_5_spec_version    = 1
pub const khr_maintenance_5_extension_name  = "VK_KHR_maintenance5"
pub type PipelineCreateFlags2KHR = u64

// Flag bits for PipelineCreateFlagBits2KHR
pub type PipelineCreateFlagBits2KHR = u64
pub const pipeline_create_2_disable_optimization_bit_khr = u64(0x00000001)
pub const pipeline_create_2_allow_derivatives_bit_khr = u64(0x00000002)
pub const pipeline_create_2_derivative_bit_khr = u64(0x00000004)
pub const pipeline_create_2_view_index_from_device_index_bit_khr = u64(0x00000008)
pub const pipeline_create_2_dispatch_base_bit_khr = u64(0x00000010)
pub const pipeline_create_2_defer_compile_bit_nv = u64(0x00000020)
pub const pipeline_create_2_capture_statistics_bit_khr = u64(0x00000040)
pub const pipeline_create_2_capture_internal_representations_bit_khr = u64(0x00000080)
pub const pipeline_create_2_fail_on_pipeline_compile_required_bit_khr = u64(0x00000100)
pub const pipeline_create_2_early_return_on_failure_bit_khr = u64(0x00000200)
pub const pipeline_create_2_link_time_optimization_bit_ext = u64(0x00000400)
pub const pipeline_create_2_retain_link_time_optimization_info_bit_ext = u64(0x00800000)
pub const pipeline_create_2_library_bit_khr = u64(0x00000800)
pub const pipeline_create_2_ray_tracing_skip_triangles_bit_khr = u64(0x00001000)
pub const pipeline_create_2_ray_tracing_skip_aabbs_bit_khr = u64(0x00002000)
pub const pipeline_create_2_ray_tracing_no_null_any_hit_shaders_bit_khr = u64(0x00004000)
pub const pipeline_create_2_ray_tracing_no_null_closest_hit_shaders_bit_khr = u64(0x00008000)
pub const pipeline_create_2_ray_tracing_no_null_miss_shaders_bit_khr = u64(0x00010000)
pub const pipeline_create_2_ray_tracing_no_null_intersection_shaders_bit_khr = u64(0x00020000)
pub const pipeline_create_2_ray_tracing_shader_group_handle_capture_replay_bit_khr = u64(0x00080000)
pub const pipeline_create_2_indirect_bindable_bit_nv = u64(0x00040000)
pub const pipeline_create_2_ray_tracing_allow_motion_bit_nv = u64(0x00100000)
pub const pipeline_create_2_rendering_fragment_shading_rate_attachment_bit_khr = u64(0x00200000)
pub const pipeline_create_2_rendering_fragment_density_map_attachment_bit_ext = u64(0x00400000)
pub const pipeline_create_2_ray_tracing_opacity_micromap_bit_ext = u64(0x01000000)
pub const pipeline_create_2_color_attachment_feedback_loop_bit_ext = u64(0x02000000)
pub const pipeline_create_2_depth_stencil_attachment_feedback_loop_bit_ext = u64(0x04000000)
pub const pipeline_create_2_no_protected_access_bit_ext = u64(0x08000000)
pub const pipeline_create_2_protected_access_only_bit_ext = u64(0x40000000)
pub const pipeline_create_2_ray_tracing_displacement_micromap_bit_nv = u64(0x10000000)
pub const pipeline_create_2_descriptor_buffer_bit_ext = u64(0x20000000)


pub type BufferUsageFlags2KHR = u64

// Flag bits for BufferUsageFlagBits2KHR
pub type BufferUsageFlagBits2KHR = u64
pub const buffer_usage_2_transfer_src_bit_khr = u64(0x00000001)
pub const buffer_usage_2_transfer_dst_bit_khr = u64(0x00000002)
pub const buffer_usage_2_uniform_texel_buffer_bit_khr = u64(0x00000004)
pub const buffer_usage_2_storage_texel_buffer_bit_khr = u64(0x00000008)
pub const buffer_usage_2_uniform_buffer_bit_khr = u64(0x00000010)
pub const buffer_usage_2_storage_buffer_bit_khr = u64(0x00000020)
pub const buffer_usage_2_index_buffer_bit_khr = u64(0x00000040)
pub const buffer_usage_2_vertex_buffer_bit_khr = u64(0x00000080)
pub const buffer_usage_2_indirect_buffer_bit_khr = u64(0x00000100)
pub const buffer_usage_2_execution_graph_scratch_bit_amdx = u64(0x02000000)
pub const buffer_usage_2_conditional_rendering_bit_ext = u64(0x00000200)
pub const buffer_usage_2_shader_binding_table_bit_khr = u64(0x00000400)
pub const buffer_usage_2_ray_tracing_bit_nv = u32(buffer_usage_2_shader_binding_table_bit_khr)
pub const buffer_usage_2_transform_feedback_buffer_bit_ext = u64(0x00000800)
pub const buffer_usage_2_transform_feedback_counter_buffer_bit_ext = u64(0x00001000)
pub const buffer_usage_2_video_decode_src_bit_khr = u64(0x00002000)
pub const buffer_usage_2_video_decode_dst_bit_khr = u64(0x00004000)
pub const buffer_usage_2_shader_device_address_bit_khr = u64(0x00020000)
pub const buffer_usage_2_acceleration_structure_build_input_read_only_bit_khr = u64(0x00080000)
pub const buffer_usage_2_acceleration_structure_storage_bit_khr = u64(0x00100000)
pub const buffer_usage_2_sampler_descriptor_buffer_bit_ext = u64(0x00200000)
pub const buffer_usage_2_resource_descriptor_buffer_bit_ext = u64(0x00400000)
pub const buffer_usage_2_push_descriptors_descriptor_buffer_bit_ext = u64(0x04000000)
pub const buffer_usage_2_micromap_build_input_read_only_bit_ext = u64(0x00800000)
pub const buffer_usage_2_micromap_storage_bit_ext = u64(0x01000000)


// PhysicalDeviceMaintenance5FeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMaintenance5FeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    maintenance5           Bool32
} 

// PhysicalDeviceMaintenance5PropertiesKHR extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceMaintenance5PropertiesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    early_fragment_multisample_coverage_after_sample_counting Bool32
    early_fragment_sample_mask_test_before_sample_counting Bool32
    depth_stencil_swizzle_one_support Bool32
    polygon_mode_point_size Bool32
    non_strict_single_pixel_wide_lines_use_parallelogram Bool32
    non_strict_wide_lines_use_parallelogram Bool32
} 

pub struct RenderingAreaInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    view_mask              u32
    color_attachment_count u32
    p_color_attachment_formats &Format
    depth_attachment_format Format
    stencil_attachment_format Format
} 

pub struct ImageSubresource2KHR {
mut:
    s_type                    StructureType
    p_next                    voidptr
    image_subresource         ImageSubresource
} 

pub struct DeviceImageSubresourceInfoKHR {
mut:
    s_type                               StructureType
    p_next                               voidptr
    p_create_info                        &ImageCreateInfo
    p_subresource                        &ImageSubresource2KHR
} 

pub struct SubresourceLayout2KHR {
mut:
    s_type                     StructureType
    p_next                     voidptr
    subresource_layout         SubresourceLayout
} 

// PipelineCreateFlags2CreateInfoKHR extends VkComputePipelineCreateInfo,VkGraphicsPipelineCreateInfo,VkRayTracingPipelineCreateInfoNV,VkRayTracingPipelineCreateInfoKHR
pub struct PipelineCreateFlags2CreateInfoKHR {
mut:
    s_type                           StructureType
    p_next                           voidptr
    flags                            PipelineCreateFlags2KHR
} 

// BufferUsageFlags2CreateInfoKHR extends VkBufferViewCreateInfo,VkBufferCreateInfo,VkPhysicalDeviceExternalBufferInfo,VkDescriptorBufferBindingInfoEXT
pub struct BufferUsageFlags2CreateInfoKHR {
mut:
    s_type                        StructureType
    p_next                        voidptr
    usage                         BufferUsageFlags2KHR
} 

type VkCmdBindIndexBuffer2KHR = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     DeviceSize,     IndexType) 

pub fn cmd_bind_index_buffer2_khr(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    size                                            DeviceSize,
    index_type                                      IndexType)  {
      f := VkCmdBindIndexBuffer2KHR((*loader_p).get_sym('vkCmdBindIndexBuffer2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindIndexBuffer2KHR': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    size,
    index_type)
}


type VkGetRenderingAreaGranularityKHR = fn (     C.Device,     &RenderingAreaInfoKHR,     &Extent2D) 

pub fn get_rendering_area_granularity_khr(
    device                                          C.Device,
    p_rendering_area_info                           &RenderingAreaInfoKHR,
    p_granularity                                   &Extent2D)  {
      f := VkGetRenderingAreaGranularityKHR((*loader_p).get_sym('vkGetRenderingAreaGranularityKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetRenderingAreaGranularityKHR': ${err}")
        return 
    })
    f(
    device,
    p_rendering_area_info,
    p_granularity)
}


type VkGetDeviceImageSubresourceLayoutKHR = fn (     C.Device,     &DeviceImageSubresourceInfoKHR,     &SubresourceLayout2KHR) 

pub fn get_device_image_subresource_layout_khr(
    device                                          C.Device,
    p_info                                          &DeviceImageSubresourceInfoKHR,
    p_layout                                        &SubresourceLayout2KHR)  {
      f := VkGetDeviceImageSubresourceLayoutKHR((*loader_p).get_sym('vkGetDeviceImageSubresourceLayoutKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceImageSubresourceLayoutKHR': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_layout)
}


type VkGetImageSubresourceLayout2KHR = fn (     C.Device,     C.Image,     &ImageSubresource2KHR,     &SubresourceLayout2KHR) 

pub fn get_image_subresource_layout2_khr(
    device                                          C.Device,
    image                                           C.Image,
    p_subresource                                   &ImageSubresource2KHR,
    p_layout                                        &SubresourceLayout2KHR)  {
      f := VkGetImageSubresourceLayout2KHR((*loader_p).get_sym('vkGetImageSubresourceLayout2KHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageSubresourceLayout2KHR': ${err}")
        return 
    })
    f(
    device,
    image,
    p_subresource,
    p_layout)
}




// VK_KHR_ray_tracing_position_fetch is a preprocessor guard. Do not pass it to API calls.
const khr_ray_tracing_position_fetch = 1
pub const khr_ray_tracing_position_fetch_spec_version = 1
pub const khr_ray_tracing_position_fetch_extension_name = "VK_KHR_ray_tracing_position_fetch"
// PhysicalDeviceRayTracingPositionFetchFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRayTracingPositionFetchFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    ray_tracing_position_fetch Bool32
} 



// VK_KHR_cooperative_matrix is a preprocessor guard. Do not pass it to API calls.
const khr_cooperative_matrix = 1
pub const khr_cooperative_matrix_spec_version = 2
pub const khr_cooperative_matrix_extension_name = "VK_KHR_cooperative_matrix"

pub enum ComponentTypeKHR {
    component_type_float16_khr = int(0)
    component_type_float32_khr = int(1)
    component_type_float64_khr = int(2)
    component_type_sint8_khr = int(3)
    component_type_sint16_khr = int(4)
    component_type_sint32_khr = int(5)
    component_type_sint64_khr = int(6)
    component_type_uint8_khr = int(7)
    component_type_uint16_khr = int(8)
    component_type_uint32_khr = int(9)
    component_type_uint64_khr = int(10)
    component_type_max_enum_khr = int(0x7FFFFFFF)
}


pub enum ScopeKHR {
    scope_device_khr = int(1)
    scope_workgroup_khr = int(2)
    scope_subgroup_khr = int(3)
    scope_queue_family_khr = int(5)
    scope_max_enum_khr = int(0x7FFFFFFF)
}

pub struct CooperativeMatrixPropertiesKHR {
mut:
    s_type                    StructureType
    p_next                    voidptr
    m_size                    u32
    n_size                    u32
    k_size                    u32
    a_type                    ComponentTypeKHR
    b_type                    ComponentTypeKHR
    c_type                    ComponentTypeKHR
    result_type               ComponentTypeKHR
    saturating_accumulation   Bool32
    scope                     ScopeKHR
} 

// PhysicalDeviceCooperativeMatrixFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceCooperativeMatrixFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    cooperative_matrix     Bool32
    cooperative_matrix_robust_buffer_access Bool32
} 

// PhysicalDeviceCooperativeMatrixPropertiesKHR extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceCooperativeMatrixPropertiesKHR {
mut:
    s_type                    StructureType
    p_next                    voidptr
    cooperative_matrix_supported_stages ShaderStageFlags
} 

type VkGetPhysicalDeviceCooperativeMatrixPropertiesKHR = fn (     C.PhysicalDevice,     &u32,     &CooperativeMatrixPropertiesKHR) Result

pub fn get_physical_device_cooperative_matrix_properties_khr(
    physical_device                                 C.PhysicalDevice,
    p_property_count                                &u32,
    p_properties                                    &CooperativeMatrixPropertiesKHR) Result {
      f := VkGetPhysicalDeviceCooperativeMatrixPropertiesKHR((*loader_p).get_sym('vkGetPhysicalDeviceCooperativeMatrixPropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceCooperativeMatrixPropertiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_property_count,
    p_properties)
}




// VK_EXT_debug_report is a preprocessor guard. Do not pass it to API calls.
const ext_debug_report = 1
pub type C.DebugReportCallbackEXT = voidptr
pub const ext_debug_report_spec_version     = 10
pub const ext_debug_report_extension_name   = "VK_EXT_debug_report"

pub enum DebugReportObjectTypeEXT {
    debug_report_object_type_unknown_ext = int(0)
    debug_report_object_type_instance_ext = int(1)
    debug_report_object_type_physical_device_ext = int(2)
    debug_report_object_type_device_ext = int(3)
    debug_report_object_type_queue_ext = int(4)
    debug_report_object_type_semaphore_ext = int(5)
    debug_report_object_type_command_buffer_ext = int(6)
    debug_report_object_type_fence_ext = int(7)
    debug_report_object_type_device_memory_ext = int(8)
    debug_report_object_type_buffer_ext = int(9)
    debug_report_object_type_image_ext = int(10)
    debug_report_object_type_event_ext = int(11)
    debug_report_object_type_query_pool_ext = int(12)
    debug_report_object_type_buffer_view_ext = int(13)
    debug_report_object_type_image_view_ext = int(14)
    debug_report_object_type_shader_module_ext = int(15)
    debug_report_object_type_pipeline_cache_ext = int(16)
    debug_report_object_type_pipeline_layout_ext = int(17)
    debug_report_object_type_render_pass_ext = int(18)
    debug_report_object_type_pipeline_ext = int(19)
    debug_report_object_type_descriptor_set_layout_ext = int(20)
    debug_report_object_type_sampler_ext = int(21)
    debug_report_object_type_descriptor_pool_ext = int(22)
    debug_report_object_type_descriptor_set_ext = int(23)
    debug_report_object_type_framebuffer_ext = int(24)
    debug_report_object_type_command_pool_ext = int(25)
    debug_report_object_type_surface_khr_ext = int(26)
    debug_report_object_type_swapchain_khr_ext = int(27)
    debug_report_object_type_debug_report_callback_ext_ext = int(28)
    debug_report_object_type_display_khr_ext = int(29)
    debug_report_object_type_display_mode_khr_ext = int(30)
    debug_report_object_type_validation_cache_ext_ext = int(33)
    debug_report_object_type_sampler_ycbcr_conversion_ext = int(1000156000)
    debug_report_object_type_descriptor_update_template_ext = int(1000085000)
    debug_report_object_type_cu_module_nvx_ext = int(1000029000)
    debug_report_object_type_cu_function_nvx_ext = int(1000029001)
    debug_report_object_type_acceleration_structure_khr_ext = int(1000150000)
    debug_report_object_type_acceleration_structure_nv_ext = int(1000165000)
    debug_report_object_type_cuda_module_nv_ext = int(1000307000)
    debug_report_object_type_cuda_function_nv_ext = int(1000307001)
    debug_report_object_type_buffer_collection_fuchsia_ext = int(1000366000)
    debug_report_object_type_max_enum_ext = int(0x7FFFFFFF)
}


pub enum DebugReportFlagBitsEXT {
    debug_report_information_bit_ext = int(0x00000001)
    debug_report_warning_bit_ext = int(0x00000002)
    debug_report_performance_warning_bit_ext = int(0x00000004)
    debug_report_error_bit_ext = int(0x00000008)
    debug_report_debug_bit_ext = int(0x00000010)
    debug_report_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type DebugReportFlagsEXT = u32
pub type PFN_vkDebugReportCallbackEXT = fn (   flags                             DebugReportFlagsEXT,   objectType                        DebugReportObjectTypeEXT,   object                            u64,   location                          usize,   messageCode                       i32,   pLayerPrefix                      &char,   pMessage                          &char,   pUserData                         voidptr) voidptr
// DebugReportCallbackCreateInfoEXT extends VkInstanceCreateInfo
pub struct DebugReportCallbackCreateInfoEXT {
mut:
    s_type                              StructureType
    p_next                              voidptr
    flags                               DebugReportFlagsEXT
    pfn_callback                        PFN_vkDebugReportCallbackEXT = unsafe { nil }
    p_user_data                         voidptr
} 

type VkCreateDebugReportCallbackEXT = fn (     C.Instance,     &DebugReportCallbackCreateInfoEXT,     &AllocationCallbacks,     &C.DebugReportCallbackEXT) Result

pub fn create_debug_report_callback_ext(
    instance                                        C.Instance,
    p_create_info                                   &DebugReportCallbackCreateInfoEXT,
    p_allocator                                     &AllocationCallbacks,
    p_callback                                      &C.DebugReportCallbackEXT) Result {
      f := VkCreateDebugReportCallbackEXT((*loader_p).get_sym('vkCreateDebugReportCallbackEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCreateDebugReportCallbackEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_callback)
}


type VkDestroyDebugReportCallbackEXT = fn (     C.Instance,     C.DebugReportCallbackEXT,     &AllocationCallbacks) 

pub fn destroy_debug_report_callback_ext(
    instance                                        C.Instance,
    callback                                        C.DebugReportCallbackEXT,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyDebugReportCallbackEXT((*loader_p).get_sym('vkDestroyDebugReportCallbackEXT'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyDebugReportCallbackEXT': ${err}")
        return 
    })
    f(
    instance,
    callback,
    p_allocator)
}


type VkDebugReportMessageEXT = fn (     C.Instance,     DebugReportFlagsEXT,     DebugReportObjectTypeEXT,     u64,     usize,     i32,     &char,     &char) 

pub fn debug_report_message_ext(
    instance                                        C.Instance,
    flags                                           DebugReportFlagsEXT,
    object_type                                     DebugReportObjectTypeEXT,
    object                                          u64,
    location                                        usize,
    message_code                                    i32,
    p_layer_prefix                                  &char,
    p_message                                       &char)  {
      f := VkDebugReportMessageEXT((*loader_p).get_sym('vkDebugReportMessageEXT'
    ) or { 
        println("Couldn't load symbol for 'vkDebugReportMessageEXT': ${err}")
        return 
    })
    f(
    instance,
    flags,
    object_type,
    object,
    location,
    message_code,
    p_layer_prefix,
    p_message)
}




// VK_NV_glsl_shader is a preprocessor guard. Do not pass it to API calls.
const nv_glsl_shader = 1
pub const nv_glsl_shader_spec_version       = 1
pub const nv_glsl_shader_extension_name     = "VK_NV_glsl_shader"


// VK_EXT_depth_range_unrestricted is a preprocessor guard. Do not pass it to API calls.
const ext_depth_range_unrestricted = 1
pub const ext_depth_range_unrestricted_spec_version = 1
pub const ext_depth_range_unrestricted_extension_name = "VK_EXT_depth_range_unrestricted"


// VK_IMG_filter_cubic is a preprocessor guard. Do not pass it to API calls.
const img_filter_cubic = 1
pub const img_filter_cubic_spec_version     = 1
pub const img_filter_cubic_extension_name   = "VK_IMG_filter_cubic"


// VK_AMD_rasterization_order is a preprocessor guard. Do not pass it to API calls.
const amd_rasterization_order = 1
pub const amd_rasterization_order_spec_version = 1
pub const amd_rasterization_order_extension_name = "VK_AMD_rasterization_order"

pub enum RasterizationOrderAMD {
    rasterization_order_strict_amd = int(0)
    rasterization_order_relaxed_amd = int(1)
    rasterization_order_max_enum_amd = int(0x7FFFFFFF)
}

// PipelineRasterizationStateRasterizationOrderAMD extends VkPipelineRasterizationStateCreateInfo
pub struct PipelineRasterizationStateRasterizationOrderAMD {
mut:
    s_type                         StructureType
    p_next                         voidptr
    rasterization_order            RasterizationOrderAMD
} 



// VK_AMD_shader_trinary_minmax is a preprocessor guard. Do not pass it to API calls.
const amd_shader_trinary_minmax = 1
pub const amd_shader_trinary_minmax_spec_version = 1
pub const amd_shader_trinary_minmax_extension_name = "VK_AMD_shader_trinary_minmax"


// VK_AMD_shader_explicit_vertex_parameter is a preprocessor guard. Do not pass it to API calls.
const amd_shader_explicit_vertex_parameter = 1
pub const amd_shader_explicit_vertex_parameter_spec_version = 1
pub const amd_shader_explicit_vertex_parameter_extension_name = "VK_AMD_shader_explicit_vertex_parameter"


// VK_EXT_debug_marker is a preprocessor guard. Do not pass it to API calls.
const ext_debug_marker = 1
pub const ext_debug_marker_spec_version     = 4
pub const ext_debug_marker_extension_name   = "VK_EXT_debug_marker"
pub struct DebugMarkerObjectNameInfoEXT {
mut:
    s_type                            StructureType
    p_next                            voidptr
    object_type                       DebugReportObjectTypeEXT
    object                            u64
    p_object_name                     &char
} 

pub struct DebugMarkerObjectTagInfoEXT {
mut:
    s_type                            StructureType
    p_next                            voidptr
    object_type                       DebugReportObjectTypeEXT
    object                            u64
    tag_name                          u64
    tag_size                          usize
    p_tag                             voidptr
} 

pub struct DebugMarkerMarkerInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    p_marker_name          &char
    color                  []f32
} 

type VkDebugMarkerSetObjectTagEXT = fn (     C.Device,     &DebugMarkerObjectTagInfoEXT) Result

pub fn debug_marker_set_object_tag_ext(
    device                                          C.Device,
    p_tag_info                                      &DebugMarkerObjectTagInfoEXT) Result {
      f := VkDebugMarkerSetObjectTagEXT((*loader_p).get_sym('vkDebugMarkerSetObjectTagEXT'
    ) or { 
        println("Couldn't load symbol for 'vkDebugMarkerSetObjectTagEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_tag_info)
}


type VkDebugMarkerSetObjectNameEXT = fn (     C.Device,     &DebugMarkerObjectNameInfoEXT) Result

pub fn debug_marker_set_object_name_ext(
    device                                          C.Device,
    p_name_info                                     &DebugMarkerObjectNameInfoEXT) Result {
      f := VkDebugMarkerSetObjectNameEXT((*loader_p).get_sym('vkDebugMarkerSetObjectNameEXT'
    ) or { 
        println("Couldn't load symbol for 'vkDebugMarkerSetObjectNameEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_name_info)
}


type VkCmdDebugMarkerBeginEXT = fn (     C.CommandBuffer,     &DebugMarkerMarkerInfoEXT) 

pub fn cmd_debug_marker_begin_ext(
    command_buffer                                  C.CommandBuffer,
    p_marker_info                                   &DebugMarkerMarkerInfoEXT)  {
      f := VkCmdDebugMarkerBeginEXT((*loader_p).get_sym('vkCmdDebugMarkerBeginEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDebugMarkerBeginEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    p_marker_info)
}


type VkCmdDebugMarkerEndEXT = fn (     C.CommandBuffer) 

pub fn cmd_debug_marker_end_ext(
    command_buffer                                  C.CommandBuffer)  {
      f := VkCmdDebugMarkerEndEXT((*loader_p).get_sym('vkCmdDebugMarkerEndEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDebugMarkerEndEXT': ${err}")
        return 
    })
    f(
    command_buffer)
}


type VkCmdDebugMarkerInsertEXT = fn (     C.CommandBuffer,     &DebugMarkerMarkerInfoEXT) 

pub fn cmd_debug_marker_insert_ext(
    command_buffer                                  C.CommandBuffer,
    p_marker_info                                   &DebugMarkerMarkerInfoEXT)  {
      f := VkCmdDebugMarkerInsertEXT((*loader_p).get_sym('vkCmdDebugMarkerInsertEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDebugMarkerInsertEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    p_marker_info)
}




// VK_AMD_gcn_shader is a preprocessor guard. Do not pass it to API calls.
const amd_gcn_shader = 1
pub const amd_gcn_shader_spec_version       = 1
pub const amd_gcn_shader_extension_name     = "VK_AMD_gcn_shader"


// VK_NV_dedicated_allocation is a preprocessor guard. Do not pass it to API calls.
const nv_dedicated_allocation = 1
pub const nv_dedicated_allocation_spec_version = 1
pub const nv_dedicated_allocation_extension_name = "VK_NV_dedicated_allocation"
// DedicatedAllocationImageCreateInfoNV extends VkImageCreateInfo
pub struct DedicatedAllocationImageCreateInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    dedicated_allocation   Bool32
} 

// DedicatedAllocationBufferCreateInfoNV extends VkBufferCreateInfo
pub struct DedicatedAllocationBufferCreateInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    dedicated_allocation   Bool32
} 

// DedicatedAllocationMemoryAllocateInfoNV extends VkMemoryAllocateInfo
pub struct DedicatedAllocationMemoryAllocateInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image                  C.Image
    buffer                 C.Buffer
} 



// VK_EXT_transform_feedback is a preprocessor guard. Do not pass it to API calls.
const ext_transform_feedback = 1
pub const ext_transform_feedback_spec_version = 1
pub const ext_transform_feedback_extension_name = "VK_EXT_transform_feedback"
pub type PipelineRasterizationStateStreamCreateFlagsEXT = u32
// PhysicalDeviceTransformFeedbackFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceTransformFeedbackFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    transform_feedback     Bool32
    geometry_streams       Bool32
} 

// PhysicalDeviceTransformFeedbackPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceTransformFeedbackPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_transform_feedback_streams u32
    max_transform_feedback_buffers u32
    max_transform_feedback_buffer_size DeviceSize
    max_transform_feedback_stream_data_size u32
    max_transform_feedback_buffer_data_size u32
    max_transform_feedback_buffer_data_stride u32
    transform_feedback_queries Bool32
    transform_feedback_streams_lines_triangles Bool32
    transform_feedback_rasterization_stream_select Bool32
    transform_feedback_draw Bool32
} 

// PipelineRasterizationStateStreamCreateInfoEXT extends VkPipelineRasterizationStateCreateInfo
pub struct PipelineRasterizationStateStreamCreateInfoEXT {
mut:
    s_type                                                  StructureType
    p_next                                                  voidptr
    flags                                                   PipelineRasterizationStateStreamCreateFlagsEXT
    rasterization_stream                                    u32
} 

type VkCmdBindTransformFeedbackBuffersEXT = fn (     C.CommandBuffer,     u32,     u32,     &C.Buffer,     &DeviceSize,     &DeviceSize) 

pub fn cmd_bind_transform_feedback_buffers_ext(
    command_buffer                                  C.CommandBuffer,
    first_binding                                   u32,
    binding_count                                   u32,
    p_buffers                                       &C.Buffer,
    p_offsets                                       &DeviceSize,
    p_sizes                                         &DeviceSize)  {
      f := VkCmdBindTransformFeedbackBuffersEXT((*loader_p).get_sym('vkCmdBindTransformFeedbackBuffersEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindTransformFeedbackBuffersEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    first_binding,
    binding_count,
    p_buffers,
    p_offsets,
    p_sizes)
}


type VkCmdBeginTransformFeedbackEXT = fn (     C.CommandBuffer,     u32,     u32,     &C.Buffer,     &DeviceSize) 

pub fn cmd_begin_transform_feedback_ext(
    command_buffer                                  C.CommandBuffer,
    first_counter_buffer                            u32,
    counter_buffer_count                            u32,
    p_counter_buffers                               &C.Buffer,
    p_counter_buffer_offsets                        &DeviceSize)  {
      f := VkCmdBeginTransformFeedbackEXT((*loader_p).get_sym('vkCmdBeginTransformFeedbackEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBeginTransformFeedbackEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    first_counter_buffer,
    counter_buffer_count,
    p_counter_buffers,
    p_counter_buffer_offsets)
}


type VkCmdEndTransformFeedbackEXT = fn (     C.CommandBuffer,     u32,     u32,     &C.Buffer,     &DeviceSize) 

pub fn cmd_end_transform_feedback_ext(
    command_buffer                                  C.CommandBuffer,
    first_counter_buffer                            u32,
    counter_buffer_count                            u32,
    p_counter_buffers                               &C.Buffer,
    p_counter_buffer_offsets                        &DeviceSize)  {
      f := VkCmdEndTransformFeedbackEXT((*loader_p).get_sym('vkCmdEndTransformFeedbackEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEndTransformFeedbackEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    first_counter_buffer,
    counter_buffer_count,
    p_counter_buffers,
    p_counter_buffer_offsets)
}


type VkCmdBeginQueryIndexedEXT = fn (     C.CommandBuffer,     C.QueryPool,     u32,     QueryControlFlags,     u32) 

pub fn cmd_begin_query_indexed_ext(
    command_buffer                                  C.CommandBuffer,
    query_pool                                      C.QueryPool,
    query                                           u32,
    flags                                           QueryControlFlags,
    index                                           u32)  {
      f := VkCmdBeginQueryIndexedEXT((*loader_p).get_sym('vkCmdBeginQueryIndexedEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBeginQueryIndexedEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    query_pool,
    query,
    flags,
    index)
}


type VkCmdEndQueryIndexedEXT = fn (     C.CommandBuffer,     C.QueryPool,     u32,     u32) 

pub fn cmd_end_query_indexed_ext(
    command_buffer                                  C.CommandBuffer,
    query_pool                                      C.QueryPool,
    query                                           u32,
    index                                           u32)  {
      f := VkCmdEndQueryIndexedEXT((*loader_p).get_sym('vkCmdEndQueryIndexedEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEndQueryIndexedEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    query_pool,
    query,
    index)
}


type VkCmdDrawIndirectByteCountEXT = fn (     C.CommandBuffer,     u32,     u32,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_indirect_byte_count_ext(
    command_buffer                                  C.CommandBuffer,
    instance_count                                  u32,
    first_instance                                  u32,
    counter_buffer                                  C.Buffer,
    counter_buffer_offset                           DeviceSize,
    counter_offset                                  u32,
    vertex_stride                                   u32)  {
      f := VkCmdDrawIndirectByteCountEXT((*loader_p).get_sym('vkCmdDrawIndirectByteCountEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawIndirectByteCountEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    instance_count,
    first_instance,
    counter_buffer,
    counter_buffer_offset,
    counter_offset,
    vertex_stride)
}




// VK_NVX_binary_import is a preprocessor guard. Do not pass it to API calls.
const nvx_binary_import = 1
pub type C.CuModuleNVX = voidptr
pub type C.CuFunctionNVX = voidptr
pub const nvx_binary_import_spec_version    = 1
pub const nvx_binary_import_extension_name  = "VK_NVX_binary_import"
pub struct CuModuleCreateInfoNVX {
mut:
    s_type                 StructureType
    p_next                 voidptr
    data_size              usize
    p_data                 voidptr
} 

pub struct CuFunctionCreateInfoNVX {
mut:
    s_type                 StructureType
    p_next                 voidptr
    vkmodule               C.CuModuleNVX
    p_name                 &char
} 

pub struct CuLaunchInfoNVX {
mut:
    s_type                     StructureType
    p_next                     voidptr
    function                   C.CuFunctionNVX
    grid_dim_x                 u32
    grid_dim_y                 u32
    grid_dim_z                 u32
    block_dim_x                u32
    block_dim_y                u32
    block_dim_z                u32
    shared_mem_bytes           u32
    param_count                usize
    p_params                   voidptr
    extra_count                usize
    p_extras                   voidptr
} 

type VkCreateCuModuleNVX = fn (     C.Device,     &CuModuleCreateInfoNVX,     &AllocationCallbacks,     &C.CuModuleNVX) Result

pub fn create_cu_module_nvx(
    device                                          C.Device,
    p_create_info                                   &CuModuleCreateInfoNVX,
    p_allocator                                     &AllocationCallbacks,
    p_module                                        &C.CuModuleNVX) Result {
      f := VkCreateCuModuleNVX((*loader_p).get_sym('vkCreateCuModuleNVX'
    ) or { 
        println("Couldn't load symbol for 'vkCreateCuModuleNVX': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_module)
}


type VkCreateCuFunctionNVX = fn (     C.Device,     &CuFunctionCreateInfoNVX,     &AllocationCallbacks,     &C.CuFunctionNVX) Result

pub fn create_cu_function_nvx(
    device                                          C.Device,
    p_create_info                                   &CuFunctionCreateInfoNVX,
    p_allocator                                     &AllocationCallbacks,
    p_function                                      &C.CuFunctionNVX) Result {
      f := VkCreateCuFunctionNVX((*loader_p).get_sym('vkCreateCuFunctionNVX'
    ) or { 
        println("Couldn't load symbol for 'vkCreateCuFunctionNVX': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_function)
}


type VkDestroyCuModuleNVX = fn (     C.Device,     C.CuModuleNVX,     &AllocationCallbacks) 

pub fn destroy_cu_module_nvx(
    device                                          C.Device,
    vkmodule                                        C.CuModuleNVX,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyCuModuleNVX((*loader_p).get_sym('vkDestroyCuModuleNVX'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyCuModuleNVX': ${err}")
        return 
    })
    f(
    device,
    vkmodule,
    p_allocator)
}


type VkDestroyCuFunctionNVX = fn (     C.Device,     C.CuFunctionNVX,     &AllocationCallbacks) 

pub fn destroy_cu_function_nvx(
    device                                          C.Device,
    function                                        C.CuFunctionNVX,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyCuFunctionNVX((*loader_p).get_sym('vkDestroyCuFunctionNVX'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyCuFunctionNVX': ${err}")
        return 
    })
    f(
    device,
    function,
    p_allocator)
}


type VkCmdCuLaunchKernelNVX = fn (     C.CommandBuffer,     &CuLaunchInfoNVX) 

pub fn cmd_cu_launch_kernel_nvx(
    command_buffer                                  C.CommandBuffer,
    p_launch_info                                   &CuLaunchInfoNVX)  {
      f := VkCmdCuLaunchKernelNVX((*loader_p).get_sym('vkCmdCuLaunchKernelNVX'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCuLaunchKernelNVX': ${err}")
        return 
    })
    f(
    command_buffer,
    p_launch_info)
}




// VK_NVX_image_view_handle is a preprocessor guard. Do not pass it to API calls.
const nvx_image_view_handle = 1
pub const nvx_image_view_handle_spec_version = 2
pub const nvx_image_view_handle_extension_name = "VK_NVX_image_view_handle"
pub struct ImageViewHandleInfoNVX {
mut:
    s_type                  StructureType
    p_next                  voidptr
    image_view              C.ImageView
    descriptor_type         DescriptorType
    sampler                 C.Sampler
} 

pub struct ImageViewAddressPropertiesNVX {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_address         DeviceAddress
    size                   DeviceSize
} 

type VkGetImageViewHandleNVX = fn (     C.Device,     &ImageViewHandleInfoNVX) u32

pub fn get_image_view_handle_nvx(
    device                                          C.Device,
    p_info                                          &ImageViewHandleInfoNVX) u32 {
      f := VkGetImageViewHandleNVX((*loader_p).get_sym("vkGetImageViewHandleNVX"
    ) or { 
        panic("Couldn't load symbol for 'vkGetImageViewHandleNVX': ${err}") })
    return f(
    device,
    p_info)
}


type VkGetImageViewAddressNVX = fn (     C.Device,     C.ImageView,     &ImageViewAddressPropertiesNVX) Result

pub fn get_image_view_address_nvx(
    device                                          C.Device,
    image_view                                      C.ImageView,
    p_properties                                    &ImageViewAddressPropertiesNVX) Result {
      f := VkGetImageViewAddressNVX((*loader_p).get_sym('vkGetImageViewAddressNVX'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageViewAddressNVX': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    image_view,
    p_properties)
}




// VK_AMD_draw_indirect_count is a preprocessor guard. Do not pass it to API calls.
const amd_draw_indirect_count = 1
pub const amd_draw_indirect_count_spec_version = 2
pub const amd_draw_indirect_count_extension_name = "VK_AMD_draw_indirect_count"
type VkCmdDrawIndirectCountAMD = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_indirect_count_amd(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    count_buffer                                    C.Buffer,
    count_buffer_offset                             DeviceSize,
    max_draw_count                                  u32,
    stride                                          u32)  {
      f := VkCmdDrawIndirectCountAMD((*loader_p).get_sym('vkCmdDrawIndirectCountAMD'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawIndirectCountAMD': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    count_buffer,
    count_buffer_offset,
    max_draw_count,
    stride)
}


type VkCmdDrawIndexedIndirectCountAMD = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_indexed_indirect_count_amd(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    count_buffer                                    C.Buffer,
    count_buffer_offset                             DeviceSize,
    max_draw_count                                  u32,
    stride                                          u32)  {
      f := VkCmdDrawIndexedIndirectCountAMD((*loader_p).get_sym('vkCmdDrawIndexedIndirectCountAMD'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawIndexedIndirectCountAMD': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    count_buffer,
    count_buffer_offset,
    max_draw_count,
    stride)
}




// VK_AMD_negative_viewport_height is a preprocessor guard. Do not pass it to API calls.
const amd_negative_viewport_height = 1
pub const amd_negative_viewport_height_spec_version = 1
pub const amd_negative_viewport_height_extension_name = "VK_AMD_negative_viewport_height"


// VK_AMD_gpu_shader_half_float is a preprocessor guard. Do not pass it to API calls.
const amd_gpu_shader_half_float = 1
pub const amd_gpu_shader_half_float_spec_version = 2
pub const amd_gpu_shader_half_float_extension_name = "VK_AMD_gpu_shader_half_float"


// VK_AMD_shader_ballot is a preprocessor guard. Do not pass it to API calls.
const amd_shader_ballot = 1
pub const amd_shader_ballot_spec_version    = 1
pub const amd_shader_ballot_extension_name  = "VK_AMD_shader_ballot"


// VK_EXT_video_encode_h264 is a preprocessor guard. Do not pass it to API calls.
const ext_video_encode_h264 = 1
pub const ext_video_encode_h264_spec_version = 12
pub const ext_video_encode_h264_extension_name = "VK_EXT_video_encode_h264"

pub enum VideoEncodeH264CapabilityFlagBitsEXT {
    video_encode_h264_capability_hrd_compliance_bit_ext = int(0x00000001)
    video_encode_h264_capability_prediction_weight_table_generated_bit_ext = int(0x00000002)
    video_encode_h264_capability_row_unaligned_slice_bit_ext = int(0x00000004)
    video_encode_h264_capability_different_slice_type_bit_ext = int(0x00000008)
    video_encode_h264_capability_b_frame_in_l0_list_bit_ext = int(0x00000010)
    video_encode_h264_capability_b_frame_in_l1_list_bit_ext = int(0x00000020)
    video_encode_h264_capability_per_picture_type_min_max_qp_bit_ext = int(0x00000040)
    video_encode_h264_capability_per_slice_constant_qp_bit_ext = int(0x00000080)
    video_encode_h264_capability_generate_prefix_nalu_bit_ext = int(0x00000100)
    video_encode_h264_capability_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type VideoEncodeH264CapabilityFlagsEXT = u32

pub enum VideoEncodeH264StdFlagBitsEXT {
    video_encode_h264_std_separate_color_plane_flag_set_bit_ext = int(0x00000001)
    video_encode_h264_std_qpprime_y_zero_transform_bypass_flag_set_bit_ext = int(0x00000002)
    video_encode_h264_std_scaling_matrix_present_flag_set_bit_ext = int(0x00000004)
    video_encode_h264_std_chroma_qp_index_offset_bit_ext = int(0x00000008)
    video_encode_h264_std_second_chroma_qp_index_offset_bit_ext = int(0x00000010)
    video_encode_h264_std_pic_init_qp_minus26_bit_ext = int(0x00000020)
    video_encode_h264_std_weighted_pred_flag_set_bit_ext = int(0x00000040)
    video_encode_h264_std_weighted_bipred_idc_explicit_bit_ext = int(0x00000080)
    video_encode_h264_std_weighted_bipred_idc_implicit_bit_ext = int(0x00000100)
    video_encode_h264_std_transform_8x8_mode_flag_set_bit_ext = int(0x00000200)
    video_encode_h264_std_direct_spatial_mv_pred_flag_unset_bit_ext = int(0x00000400)
    video_encode_h264_std_entropy_coding_mode_flag_unset_bit_ext = int(0x00000800)
    video_encode_h264_std_entropy_coding_mode_flag_set_bit_ext = int(0x00001000)
    video_encode_h264_std_direct_8x8_inference_flag_unset_bit_ext = int(0x00002000)
    video_encode_h264_std_constrained_intra_pred_flag_set_bit_ext = int(0x00004000)
    video_encode_h264_std_deblocking_filter_disabled_bit_ext = int(0x00008000)
    video_encode_h264_std_deblocking_filter_enabled_bit_ext = int(0x00010000)
    video_encode_h264_std_deblocking_filter_partial_bit_ext = int(0x00020000)
    video_encode_h264_std_slice_qp_delta_bit_ext = int(0x00080000)
    video_encode_h264_std_different_slice_qp_delta_bit_ext = int(0x00100000)
    video_encode_h264_std_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type VideoEncodeH264StdFlagsEXT = u32

pub enum VideoEncodeH264RateControlFlagBitsEXT {
    video_encode_h264_rate_control_attempt_hrd_compliance_bit_ext = int(0x00000001)
    video_encode_h264_rate_control_regular_gop_bit_ext = int(0x00000002)
    video_encode_h264_rate_control_reference_pattern_flat_bit_ext = int(0x00000004)
    video_encode_h264_rate_control_reference_pattern_dyadic_bit_ext = int(0x00000008)
    video_encode_h264_rate_control_temporal_layer_pattern_dyadic_bit_ext = int(0x00000010)
    video_encode_h264_rate_control_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type VideoEncodeH264RateControlFlagsEXT = u32
// VideoEncodeH264CapabilitiesEXT extends VkVideoCapabilitiesKHR
pub struct VideoEncodeH264CapabilitiesEXT {
mut:
    s_type                                     StructureType
    p_next                                     voidptr
    flags                                      VideoEncodeH264CapabilityFlagsEXT
    max_level_idc                              C.StdVideoH264LevelIdc
    max_slice_count                            u32
    max_p_picture_l0_reference_count           u32
    max_b_picture_l0_reference_count           u32
    max_l1_reference_count                     u32
    max_temporal_layer_count                   u32
    expect_dyadic_temporal_layer_pattern       Bool32
    min_qp                                     i32
    max_qp                                     i32
    prefers_gop_remaining_frames               Bool32
    requires_gop_remaining_frames              Bool32
    std_syntax_flags                           VideoEncodeH264StdFlagsEXT
} 

pub struct VideoEncodeH264QpEXT {
mut:
    qp_i           i32
    qp_p           i32
    qp_b           i32
} 

// VideoEncodeH264QualityLevelPropertiesEXT extends VkVideoEncodeQualityLevelPropertiesKHR
pub struct VideoEncodeH264QualityLevelPropertiesEXT {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    preferred_rate_control_flags                VideoEncodeH264RateControlFlagsEXT
    preferred_gop_frame_count                   u32
    preferred_idr_period                        u32
    preferred_consecutive_b_frame_count         u32
    preferred_temporal_layer_count              u32
    preferred_constant_qp                       VideoEncodeH264QpEXT
    preferred_max_l0_reference_count            u32
    preferred_max_l1_reference_count            u32
    preferred_std_entropy_coding_mode_flag      Bool32
} 

// VideoEncodeH264SessionCreateInfoEXT extends VkVideoSessionCreateInfoKHR
pub struct VideoEncodeH264SessionCreateInfoEXT {
mut:
    s_type                      StructureType
    p_next                      voidptr
    use_max_level_idc           Bool32
    max_level_idc               C.StdVideoH264LevelIdc
} 

// VideoEncodeH264SessionParametersAddInfoEXT extends VkVideoSessionParametersUpdateInfoKHR
pub struct VideoEncodeH264SessionParametersAddInfoEXT {
mut:
    s_type                                         StructureType
    p_next                                         voidptr
    std_sps_count                                  u32
    p_std_sp_ss                                    &C.StdVideoH264SequenceParameterSet
    std_pps_count                                  u32
    p_std_pp_ss                                    &C.StdVideoH264PictureParameterSet
} 

// VideoEncodeH264SessionParametersCreateInfoEXT extends VkVideoSessionParametersCreateInfoKHR
pub struct VideoEncodeH264SessionParametersCreateInfoEXT {
mut:
    s_type                                                     StructureType
    p_next                                                     voidptr
    max_std_sps_count                                          u32
    max_std_pps_count                                          u32
    p_parameters_add_info                                      &VideoEncodeH264SessionParametersAddInfoEXT
} 

// VideoEncodeH264SessionParametersGetInfoEXT extends VkVideoEncodeSessionParametersGetInfoKHR
pub struct VideoEncodeH264SessionParametersGetInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    write_std_sps          Bool32
    write_std_pps          Bool32
    std_sps_id             u32
    std_pps_id             u32
} 

// VideoEncodeH264SessionParametersFeedbackInfoEXT extends VkVideoEncodeSessionParametersFeedbackInfoKHR
pub struct VideoEncodeH264SessionParametersFeedbackInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    has_std_sps_overrides  Bool32
    has_std_pps_overrides  Bool32
} 

pub struct VideoEncodeH264NaluSliceInfoEXT {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    constant_qp                                 i32
    p_std_slice_header                          &C.StdVideoEncodeH264SliceHeader
} 

// VideoEncodeH264PictureInfoEXT extends VkVideoEncodeInfoKHR
pub struct VideoEncodeH264PictureInfoEXT {
mut:
    s_type                                          StructureType
    p_next                                          voidptr
    nalu_slice_entry_count                          u32
    p_nalu_slice_entries                            &VideoEncodeH264NaluSliceInfoEXT
    p_std_picture_info                              &C.StdVideoEncodeH264PictureInfo
    generate_prefix_nalu                            Bool32
} 

// VideoEncodeH264DpbSlotInfoEXT extends VkVideoReferenceSlotInfoKHR
pub struct VideoEncodeH264DpbSlotInfoEXT {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    p_std_reference_info                          &C.StdVideoEncodeH264ReferenceInfo
} 

// VideoEncodeH264ProfileInfoEXT extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub struct VideoEncodeH264ProfileInfoEXT {
mut:
    s_type                        StructureType
    p_next                        voidptr
    std_profile_idc               C.StdVideoH264ProfileIdc
} 

// VideoEncodeH264RateControlInfoEXT extends VkVideoCodingControlInfoKHR,VkVideoBeginCodingInfoKHR
pub struct VideoEncodeH264RateControlInfoEXT {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    flags                                       VideoEncodeH264RateControlFlagsEXT
    gop_frame_count                             u32
    idr_period                                  u32
    consecutive_b_frame_count                   u32
    temporal_layer_count                        u32
} 

pub struct VideoEncodeH264FrameSizeEXT {
mut:
    frame_i_size    u32
    frame_p_size    u32
    frame_b_size    u32
} 

// VideoEncodeH264RateControlLayerInfoEXT extends VkVideoEncodeRateControlLayerInfoKHR
pub struct VideoEncodeH264RateControlLayerInfoEXT {
mut:
    s_type                               StructureType
    p_next                               voidptr
    use_min_qp                           Bool32
    min_qp                               VideoEncodeH264QpEXT
    use_max_qp                           Bool32
    max_qp                               VideoEncodeH264QpEXT
    use_max_frame_size                   Bool32
    max_frame_size                       VideoEncodeH264FrameSizeEXT
} 

// VideoEncodeH264GopRemainingFrameInfoEXT extends VkVideoBeginCodingInfoKHR
pub struct VideoEncodeH264GopRemainingFrameInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    use_gop_remaining_frames Bool32
    gop_remaining_i        u32
    gop_remaining_p        u32
    gop_remaining_b        u32
} 



// VK_EXT_video_encode_h265 is a preprocessor guard. Do not pass it to API calls.
const ext_video_encode_h265 = 1
pub const ext_video_encode_h265_spec_version = 12
pub const ext_video_encode_h265_extension_name = "VK_EXT_video_encode_h265"

pub enum VideoEncodeH265CapabilityFlagBitsEXT {
    video_encode_h265_capability_hrd_compliance_bit_ext = int(0x00000001)
    video_encode_h265_capability_prediction_weight_table_generated_bit_ext = int(0x00000002)
    video_encode_h265_capability_row_unaligned_slice_segment_bit_ext = int(0x00000004)
    video_encode_h265_capability_different_slice_segment_type_bit_ext = int(0x00000008)
    video_encode_h265_capability_b_frame_in_l0_list_bit_ext = int(0x00000010)
    video_encode_h265_capability_b_frame_in_l1_list_bit_ext = int(0x00000020)
    video_encode_h265_capability_per_picture_type_min_max_qp_bit_ext = int(0x00000040)
    video_encode_h265_capability_per_slice_segment_constant_qp_bit_ext = int(0x00000080)
    video_encode_h265_capability_multiple_tiles_per_slice_segment_bit_ext = int(0x00000100)
    video_encode_h265_capability_multiple_slice_segments_per_tile_bit_ext = int(0x00000200)
    video_encode_h265_capability_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type VideoEncodeH265CapabilityFlagsEXT = u32

pub enum VideoEncodeH265StdFlagBitsEXT {
    video_encode_h265_std_separate_color_plane_flag_set_bit_ext = int(0x00000001)
    video_encode_h265_std_sample_adaptive_offset_enabled_flag_set_bit_ext = int(0x00000002)
    video_encode_h265_std_scaling_list_data_present_flag_set_bit_ext = int(0x00000004)
    video_encode_h265_std_pcm_enabled_flag_set_bit_ext = int(0x00000008)
    video_encode_h265_std_sps_temporal_mvp_enabled_flag_set_bit_ext = int(0x00000010)
    video_encode_h265_std_init_qp_minus26_bit_ext = int(0x00000020)
    video_encode_h265_std_weighted_pred_flag_set_bit_ext = int(0x00000040)
    video_encode_h265_std_weighted_bipred_flag_set_bit_ext = int(0x00000080)
    video_encode_h265_std_log2_parallel_merge_level_minus2_bit_ext = int(0x00000100)
    video_encode_h265_std_sign_data_hiding_enabled_flag_set_bit_ext = int(0x00000200)
    video_encode_h265_std_transform_skip_enabled_flag_set_bit_ext = int(0x00000400)
    video_encode_h265_std_transform_skip_enabled_flag_unset_bit_ext = int(0x00000800)
    video_encode_h265_std_pps_slice_chroma_qp_offsets_present_flag_set_bit_ext = int(0x00001000)
    video_encode_h265_std_transquant_bypass_enabled_flag_set_bit_ext = int(0x00002000)
    video_encode_h265_std_constrained_intra_pred_flag_set_bit_ext = int(0x00004000)
    video_encode_h265_std_entropy_coding_sync_enabled_flag_set_bit_ext = int(0x00008000)
    video_encode_h265_std_deblocking_filter_override_enabled_flag_set_bit_ext = int(0x00010000)
    video_encode_h265_std_dependent_slice_segments_enabled_flag_set_bit_ext = int(0x00020000)
    video_encode_h265_std_dependent_slice_segment_flag_set_bit_ext = int(0x00040000)
    video_encode_h265_std_slice_qp_delta_bit_ext = int(0x00080000)
    video_encode_h265_std_different_slice_qp_delta_bit_ext = int(0x00100000)
    video_encode_h265_std_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type VideoEncodeH265StdFlagsEXT = u32

pub enum VideoEncodeH265CtbSizeFlagBitsEXT {
    video_encode_h265_ctb_size_16_bit_ext = int(0x00000001)
    video_encode_h265_ctb_size_32_bit_ext = int(0x00000002)
    video_encode_h265_ctb_size_64_bit_ext = int(0x00000004)
    video_encode_h265_ctb_size_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type VideoEncodeH265CtbSizeFlagsEXT = u32

pub enum VideoEncodeH265TransformBlockSizeFlagBitsEXT {
    video_encode_h265_transform_block_size_4_bit_ext = int(0x00000001)
    video_encode_h265_transform_block_size_8_bit_ext = int(0x00000002)
    video_encode_h265_transform_block_size_16_bit_ext = int(0x00000004)
    video_encode_h265_transform_block_size_32_bit_ext = int(0x00000008)
    video_encode_h265_transform_block_size_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type VideoEncodeH265TransformBlockSizeFlagsEXT = u32

pub enum VideoEncodeH265RateControlFlagBitsEXT {
    video_encode_h265_rate_control_attempt_hrd_compliance_bit_ext = int(0x00000001)
    video_encode_h265_rate_control_regular_gop_bit_ext = int(0x00000002)
    video_encode_h265_rate_control_reference_pattern_flat_bit_ext = int(0x00000004)
    video_encode_h265_rate_control_reference_pattern_dyadic_bit_ext = int(0x00000008)
    video_encode_h265_rate_control_temporal_sub_layer_pattern_dyadic_bit_ext = int(0x00000010)
    video_encode_h265_rate_control_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type VideoEncodeH265RateControlFlagsEXT = u32
// VideoEncodeH265CapabilitiesEXT extends VkVideoCapabilitiesKHR
pub struct VideoEncodeH265CapabilitiesEXT {
mut:
    s_type                                             StructureType
    p_next                                             voidptr
    flags                                              VideoEncodeH265CapabilityFlagsEXT
    max_level_idc                                      u32
    max_slice_segment_count                            u32
    max_tiles                                          Extent2D
    ctb_sizes                                          VideoEncodeH265CtbSizeFlagsEXT
    transform_block_sizes                              VideoEncodeH265TransformBlockSizeFlagsEXT
    max_p_picture_l0_reference_count                   u32
    max_b_picture_l0_reference_count                   u32
    max_l1_reference_count                             u32
    max_sub_layer_count                                u32
    expect_dyadic_temporal_sub_layer_pattern           Bool32
    min_qp                                             i32
    max_qp                                             i32
    prefers_gop_remaining_frames                       Bool32
    requires_gop_remaining_frames                      Bool32
    std_syntax_flags                                   VideoEncodeH265StdFlagsEXT
} 

// VideoEncodeH265SessionCreateInfoEXT extends VkVideoSessionCreateInfoKHR
pub struct VideoEncodeH265SessionCreateInfoEXT {
mut:
    s_type                      StructureType
    p_next                      voidptr
    use_max_level_idc           Bool32
    max_level_idc               u32
} 

pub struct VideoEncodeH265QpEXT {
mut:
    qp_i           i32
    qp_p           i32
    qp_b           i32
} 

// VideoEncodeH265QualityLevelPropertiesEXT extends VkVideoEncodeQualityLevelPropertiesKHR
pub struct VideoEncodeH265QualityLevelPropertiesEXT {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    preferred_rate_control_flags                VideoEncodeH265RateControlFlagsEXT
    preferred_gop_frame_count                   u32
    preferred_idr_period                        u32
    preferred_consecutive_b_frame_count         u32
    preferred_sub_layer_count                   u32
    preferred_constant_qp                       VideoEncodeH265QpEXT
    preferred_max_l0_reference_count            u32
    preferred_max_l1_reference_count            u32
} 

// VideoEncodeH265SessionParametersAddInfoEXT extends VkVideoSessionParametersUpdateInfoKHR
pub struct VideoEncodeH265SessionParametersAddInfoEXT {
mut:
    s_type                                         StructureType
    p_next                                         voidptr
    std_vps_count                                  u32
    p_std_vp_ss                                    &C.StdVideoH265VideoParameterSet
    std_sps_count                                  u32
    p_std_sp_ss                                    &C.StdVideoH265SequenceParameterSet
    std_pps_count                                  u32
    p_std_pp_ss                                    &C.StdVideoH265PictureParameterSet
} 

// VideoEncodeH265SessionParametersCreateInfoEXT extends VkVideoSessionParametersCreateInfoKHR
pub struct VideoEncodeH265SessionParametersCreateInfoEXT {
mut:
    s_type                                                     StructureType
    p_next                                                     voidptr
    max_std_vps_count                                          u32
    max_std_sps_count                                          u32
    max_std_pps_count                                          u32
    p_parameters_add_info                                      &VideoEncodeH265SessionParametersAddInfoEXT
} 

// VideoEncodeH265SessionParametersGetInfoEXT extends VkVideoEncodeSessionParametersGetInfoKHR
pub struct VideoEncodeH265SessionParametersGetInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    write_std_vps          Bool32
    write_std_sps          Bool32
    write_std_pps          Bool32
    std_vps_id             u32
    std_sps_id             u32
    std_pps_id             u32
} 

// VideoEncodeH265SessionParametersFeedbackInfoEXT extends VkVideoEncodeSessionParametersFeedbackInfoKHR
pub struct VideoEncodeH265SessionParametersFeedbackInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    has_std_vps_overrides  Bool32
    has_std_sps_overrides  Bool32
    has_std_pps_overrides  Bool32
} 

pub struct VideoEncodeH265NaluSliceSegmentInfoEXT {
mut:
    s_type                                             StructureType
    p_next                                             voidptr
    constant_qp                                        i32
    p_std_slice_segment_header                         &C.StdVideoEncodeH265SliceSegmentHeader
} 

// VideoEncodeH265PictureInfoEXT extends VkVideoEncodeInfoKHR
pub struct VideoEncodeH265PictureInfoEXT {
mut:
    s_type                                                 StructureType
    p_next                                                 voidptr
    nalu_slice_segment_entry_count                         u32
    p_nalu_slice_segment_entries                           &VideoEncodeH265NaluSliceSegmentInfoEXT
    p_std_picture_info                                     &C.StdVideoEncodeH265PictureInfo
} 

// VideoEncodeH265DpbSlotInfoEXT extends VkVideoReferenceSlotInfoKHR
pub struct VideoEncodeH265DpbSlotInfoEXT {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    p_std_reference_info                          &C.StdVideoEncodeH265ReferenceInfo
} 

// VideoEncodeH265ProfileInfoEXT extends VkVideoProfileInfoKHR,VkQueryPoolCreateInfo
pub struct VideoEncodeH265ProfileInfoEXT {
mut:
    s_type                        StructureType
    p_next                        voidptr
    std_profile_idc               C.StdVideoH265ProfileIdc
} 

// VideoEncodeH265RateControlInfoEXT extends VkVideoCodingControlInfoKHR,VkVideoBeginCodingInfoKHR
pub struct VideoEncodeH265RateControlInfoEXT {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    flags                                       VideoEncodeH265RateControlFlagsEXT
    gop_frame_count                             u32
    idr_period                                  u32
    consecutive_b_frame_count                   u32
    sub_layer_count                             u32
} 

pub struct VideoEncodeH265FrameSizeEXT {
mut:
    frame_i_size    u32
    frame_p_size    u32
    frame_b_size    u32
} 

// VideoEncodeH265RateControlLayerInfoEXT extends VkVideoEncodeRateControlLayerInfoKHR
pub struct VideoEncodeH265RateControlLayerInfoEXT {
mut:
    s_type                               StructureType
    p_next                               voidptr
    use_min_qp                           Bool32
    min_qp                               VideoEncodeH265QpEXT
    use_max_qp                           Bool32
    max_qp                               VideoEncodeH265QpEXT
    use_max_frame_size                   Bool32
    max_frame_size                       VideoEncodeH265FrameSizeEXT
} 

// VideoEncodeH265GopRemainingFrameInfoEXT extends VkVideoBeginCodingInfoKHR
pub struct VideoEncodeH265GopRemainingFrameInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    use_gop_remaining_frames Bool32
    gop_remaining_i        u32
    gop_remaining_p        u32
    gop_remaining_b        u32
} 



// VK_AMD_texture_gather_bias_lod is a preprocessor guard. Do not pass it to API calls.
const amd_texture_gather_bias_lod = 1
pub const amd_texture_gather_bias_lod_spec_version = 1
pub const amd_texture_gather_bias_lod_extension_name = "VK_AMD_texture_gather_bias_lod"
// TextureLODGatherFormatPropertiesAMD extends VkImageFormatProperties2
pub struct TextureLODGatherFormatPropertiesAMD {
mut:
    s_type                 StructureType
    p_next                 voidptr
    supports_texture_gather_lod_bias_amd Bool32
} 



// VK_AMD_shader_info is a preprocessor guard. Do not pass it to API calls.
const amd_shader_info = 1
pub const amd_shader_info_spec_version      = 1
pub const amd_shader_info_extension_name    = "VK_AMD_shader_info"

pub enum ShaderInfoTypeAMD {
    shader_info_type_statistics_amd = int(0)
    shader_info_type_binary_amd = int(1)
    shader_info_type_disassembly_amd = int(2)
    shader_info_type_max_enum_amd = int(0x7FFFFFFF)
}

pub struct ShaderResourceUsageAMD {
mut:
    num_used_vgprs  u32
    num_used_sgprs  u32
    lds_size_per_local_work_group u32
    lds_usage_size_in_bytes usize
    scratch_mem_usage_in_bytes usize
} 

pub struct ShaderStatisticsInfoAMD {
mut:
    shader_stage_mask               ShaderStageFlags
    resource_usage                  ShaderResourceUsageAMD
    num_physical_vgprs              u32
    num_physical_sgprs              u32
    num_available_vgprs             u32
    num_available_sgprs             u32
    compute_work_group_size         []u32
} 

type VkGetShaderInfoAMD = fn (     C.Device,     C.Pipeline,     ShaderStageFlagBits,     ShaderInfoTypeAMD,     &usize,     voidptr) Result

pub fn get_shader_info_amd(
    device                                          C.Device,
    pipeline                                        C.Pipeline,
    shader_stage                                    ShaderStageFlagBits,
    info_type                                       ShaderInfoTypeAMD,
    p_info_size                                     &usize,
    p_info                                          voidptr) Result {
      f := VkGetShaderInfoAMD((*loader_p).get_sym('vkGetShaderInfoAMD'
    ) or { 
        println("Couldn't load symbol for 'vkGetShaderInfoAMD': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    pipeline,
    shader_stage,
    info_type,
    p_info_size,
    p_info)
}




// VK_AMD_shader_image_load_store_lod is a preprocessor guard. Do not pass it to API calls.
const amd_shader_image_load_store_lod = 1
pub const amd_shader_image_load_store_lod_spec_version = 1
pub const amd_shader_image_load_store_lod_extension_name = "VK_AMD_shader_image_load_store_lod"


// VK_GGP_stream_descriptor_surface is a preprocessor guard. Do not pass it to API calls.
const ggp_stream_descriptor_surface = 1
pub const ggp_stream_descriptor_surface_spec_version = 1
pub const ggp_stream_descriptor_surface_extension_name = "VK_GGP_stream_descriptor_surface"
pub type StreamDescriptorSurfaceCreateFlagsGGP = u32
pub struct StreamDescriptorSurfaceCreateInfoGGP {
mut:
    s_type                                         StructureType
    p_next                                         voidptr
    flags                                          StreamDescriptorSurfaceCreateFlagsGGP
    stream_descriptor                              voidptr
} 

type VkCreateStreamDescriptorSurfaceGGP = fn (     C.Instance,     &StreamDescriptorSurfaceCreateInfoGGP,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_stream_descriptor_surface_ggp(
    instance                                        C.Instance,
    p_create_info                                   &StreamDescriptorSurfaceCreateInfoGGP,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateStreamDescriptorSurfaceGGP((*loader_p).get_sym('vkCreateStreamDescriptorSurfaceGGP'
    ) or { 
        println("Couldn't load symbol for 'vkCreateStreamDescriptorSurfaceGGP': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}




// VK_NV_corner_sampled_image is a preprocessor guard. Do not pass it to API calls.
const nv_corner_sampled_image = 1
pub const nv_corner_sampled_image_spec_version = 2
pub const nv_corner_sampled_image_extension_name = "VK_NV_corner_sampled_image"
// PhysicalDeviceCornerSampledImageFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceCornerSampledImageFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    corner_sampled_image   Bool32
} 



// VK_IMG_format_pvrtc is a preprocessor guard. Do not pass it to API calls.
const img_format_pvrtc = 1
pub const img_format_pvrtc_spec_version     = 1
pub const img_format_pvrtc_extension_name   = "VK_IMG_format_pvrtc"


// VK_NV_external_memory_capabilities is a preprocessor guard. Do not pass it to API calls.
const nv_external_memory_capabilities = 1
pub const nv_external_memory_capabilities_spec_version = 1
pub const nv_external_memory_capabilities_extension_name = "VK_NV_external_memory_capabilities"

pub enum ExternalMemoryHandleTypeFlagBitsNV {
    external_memory_handle_type_opaque_win32_bit_nv = int(0x00000001)
    external_memory_handle_type_opaque_win32_kmt_bit_nv = int(0x00000002)
    external_memory_handle_type_d3d11_image_bit_nv = int(0x00000004)
    external_memory_handle_type_d3d11_image_kmt_bit_nv = int(0x00000008)
    external_memory_handle_type_flag_bits_max_enum_nv = int(0x7FFFFFFF)
}

pub type ExternalMemoryHandleTypeFlagsNV = u32

pub enum ExternalMemoryFeatureFlagBitsNV {
    external_memory_feature_dedicated_only_bit_nv = int(0x00000001)
    external_memory_feature_exportable_bit_nv = int(0x00000002)
    external_memory_feature_importable_bit_nv = int(0x00000004)
    external_memory_feature_flag_bits_max_enum_nv = int(0x7FFFFFFF)
}

pub type ExternalMemoryFeatureFlagsNV = u32
pub struct ExternalImageFormatPropertiesNV {
mut:
    image_format_properties                  ImageFormatProperties
    external_memory_features                 ExternalMemoryFeatureFlagsNV
    export_from_imported_handle_types        ExternalMemoryHandleTypeFlagsNV
    compatible_handle_types                  ExternalMemoryHandleTypeFlagsNV
} 

type VkGetPhysicalDeviceExternalImageFormatPropertiesNV = fn (     C.PhysicalDevice,     Format,     ImageType,     ImageTiling,     ImageUsageFlags,     ImageCreateFlags,     ExternalMemoryHandleTypeFlagsNV,     &ExternalImageFormatPropertiesNV) Result

pub fn get_physical_device_external_image_format_properties_nv(
    physical_device                                 C.PhysicalDevice,
    format                                          Format,
    vktype                                          ImageType,
    tiling                                          ImageTiling,
    usage                                           ImageUsageFlags,
    flags                                           ImageCreateFlags,
    external_handle_type                            ExternalMemoryHandleTypeFlagsNV,
    p_external_image_format_properties              &ExternalImageFormatPropertiesNV) Result {
      f := VkGetPhysicalDeviceExternalImageFormatPropertiesNV((*loader_p).get_sym('vkGetPhysicalDeviceExternalImageFormatPropertiesNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceExternalImageFormatPropertiesNV': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    format,
    vktype,
    tiling,
    usage,
    flags,
    external_handle_type,
    p_external_image_format_properties)
}




// VK_NV_external_memory is a preprocessor guard. Do not pass it to API calls.
const nv_external_memory = 1
pub const nv_external_memory_spec_version   = 1
pub const nv_external_memory_extension_name = "VK_NV_external_memory"
// ExternalMemoryImageCreateInfoNV extends VkImageCreateInfo
pub struct ExternalMemoryImageCreateInfoNV {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    handle_types                             ExternalMemoryHandleTypeFlagsNV
} 

// ExportMemoryAllocateInfoNV extends VkMemoryAllocateInfo
pub struct ExportMemoryAllocateInfoNV {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    handle_types                             ExternalMemoryHandleTypeFlagsNV
} 



// VK_NV_external_memory_win32 is a preprocessor guard. Do not pass it to API calls.
const nv_external_memory_win32 = 1
pub const nv_external_memory_win32_spec_version = 1
pub const nv_external_memory_win32_extension_name = "VK_NV_external_memory_win32"
// ImportMemoryWin32HandleInfoNV extends VkMemoryAllocateInfo
pub struct ImportMemoryWin32HandleInfoNV {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    handle_type                              ExternalMemoryHandleTypeFlagsNV
    handle                                   voidptr
} 

// ExportMemoryWin32HandleInfoNV extends VkMemoryAllocateInfo
pub struct ExportMemoryWin32HandleInfoNV {
mut:
    s_type                            StructureType
    p_next                            voidptr
    p_attributes                      voidptr
    dw_access                         u32
} 

type VkGetMemoryWin32HandleNV = fn (     C.Device,     C.DeviceMemory,     ExternalMemoryHandleTypeFlagsNV,     &voidptr) Result

pub fn get_memory_win32_handle_nv(
    device                                          C.Device,
    memory                                          C.DeviceMemory,
    handle_type                                     ExternalMemoryHandleTypeFlagsNV,
    p_handle                                        &voidptr) Result {
      f := VkGetMemoryWin32HandleNV((*loader_p).get_sym('vkGetMemoryWin32HandleNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetMemoryWin32HandleNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    memory,
    handle_type,
    p_handle)
}




// VK_NV_win32_keyed_mutex is a preprocessor guard. Do not pass it to API calls.
const nv_win32_keyed_mutex = 1
pub const nv_win32_keyed_mutex_spec_version = 2
pub const nv_win32_keyed_mutex_extension_name = "VK_NV_win32_keyed_mutex"
// Win32KeyedMutexAcquireReleaseInfoNV extends VkSubmitInfo,VkSubmitInfo2
pub struct Win32KeyedMutexAcquireReleaseInfoNV {
mut:
    s_type                       StructureType
    p_next                       voidptr
    acquire_count                u32
    p_acquire_syncs              &C.DeviceMemory
    p_acquire_keys               &u64
    p_acquire_timeout_milliseconds &u32
    release_count                u32
    p_release_syncs              &C.DeviceMemory
    p_release_keys               &u64
} 



// VK_EXT_validation_flags is a preprocessor guard. Do not pass it to API calls.
const ext_validation_flags = 1
pub const ext_validation_flags_spec_version = 3
pub const ext_validation_flags_extension_name = "VK_EXT_validation_flags"

pub enum ValidationCheckEXT {
    validation_check_all_ext = int(0)
    validation_check_shaders_ext = int(1)
    validation_check_max_enum_ext = int(0x7FFFFFFF)
}

// ValidationFlagsEXT extends VkInstanceCreateInfo
pub struct ValidationFlagsEXT {
mut:
    s_type                             StructureType
    p_next                             voidptr
    disabled_validation_check_count    u32
    p_disabled_validation_checks       &ValidationCheckEXT
} 



// VK_NN_vi_surface is a preprocessor guard. Do not pass it to API calls.
const nn_vi_surface = 1
pub const nn_vi_surface_spec_version        = 1
pub const nn_vi_surface_extension_name      = "VK_NN_vi_surface"
pub type ViSurfaceCreateFlagsNN = u32
pub struct ViSurfaceCreateInfoNN {
mut:
    s_type                          StructureType
    p_next                          voidptr
    flags                           ViSurfaceCreateFlagsNN
    window                          voidptr
} 

type VkCreateViSurfaceNN = fn (     C.Instance,     &ViSurfaceCreateInfoNN,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_vi_surface_nn(
    instance                                        C.Instance,
    p_create_info                                   &ViSurfaceCreateInfoNN,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateViSurfaceNN((*loader_p).get_sym('vkCreateViSurfaceNN'
    ) or { 
        println("Couldn't load symbol for 'vkCreateViSurfaceNN': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}




// VK_EXT_shader_subgroup_ballot is a preprocessor guard. Do not pass it to API calls.
const ext_shader_subgroup_ballot = 1
pub const ext_shader_subgroup_ballot_spec_version = 1
pub const ext_shader_subgroup_ballot_extension_name = "VK_EXT_shader_subgroup_ballot"


// VK_EXT_shader_subgroup_vote is a preprocessor guard. Do not pass it to API calls.
const ext_shader_subgroup_vote = 1
pub const ext_shader_subgroup_vote_spec_version = 1
pub const ext_shader_subgroup_vote_extension_name = "VK_EXT_shader_subgroup_vote"


// VK_EXT_texture_compression_astc_hdr is a preprocessor guard. Do not pass it to API calls.
const ext_texture_compression_astc_hdr = 1
pub const ext_texture_compression_astc_hdr_spec_version = 1
pub const ext_texture_compression_astc_hdr_extension_name = "VK_EXT_texture_compression_astc_hdr"
pub type PhysicalDeviceTextureCompressionASTCHDRFeaturesEXT = PhysicalDeviceTextureCompressionASTCHDRFeatures



// VK_EXT_astc_decode_mode is a preprocessor guard. Do not pass it to API calls.
const ext_astc_decode_mode = 1
pub const ext_astc_decode_mode_spec_version = 1
pub const ext_astc_decode_mode_extension_name = "VK_EXT_astc_decode_mode"
// ImageViewASTCDecodeModeEXT extends VkImageViewCreateInfo
pub struct ImageViewASTCDecodeModeEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    decode_mode            Format
} 

// PhysicalDeviceASTCDecodeFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceASTCDecodeFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    decode_mode_shared_exponent Bool32
} 



// VK_EXT_pipeline_robustness is a preprocessor guard. Do not pass it to API calls.
const ext_pipeline_robustness = 1
pub const ext_pipeline_robustness_spec_version = 1
pub const ext_pipeline_robustness_extension_name = "VK_EXT_pipeline_robustness"

pub enum PipelineRobustnessBufferBehaviorEXT {
    pipeline_robustness_buffer_behavior_device_default_ext = int(0)
    pipeline_robustness_buffer_behavior_disabled_ext = int(1)
    pipeline_robustness_buffer_behavior_robust_buffer_access_ext = int(2)
    pipeline_robustness_buffer_behavior_robust_buffer_access_2_ext = int(3)
    pipeline_robustness_buffer_behavior_max_enum_ext = int(0x7FFFFFFF)
}


pub enum PipelineRobustnessImageBehaviorEXT {
    pipeline_robustness_image_behavior_device_default_ext = int(0)
    pipeline_robustness_image_behavior_disabled_ext = int(1)
    pipeline_robustness_image_behavior_robust_image_access_ext = int(2)
    pipeline_robustness_image_behavior_robust_image_access_2_ext = int(3)
    pipeline_robustness_image_behavior_max_enum_ext = int(0x7FFFFFFF)
}

// PhysicalDevicePipelineRobustnessFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePipelineRobustnessFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pipeline_robustness    Bool32
} 

// PhysicalDevicePipelineRobustnessPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDevicePipelineRobustnessPropertiesEXT {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    default_robustness_storage_buffers           PipelineRobustnessBufferBehaviorEXT
    default_robustness_uniform_buffers           PipelineRobustnessBufferBehaviorEXT
    default_robustness_vertex_inputs             PipelineRobustnessBufferBehaviorEXT
    default_robustness_images                    PipelineRobustnessImageBehaviorEXT
} 

// PipelineRobustnessCreateInfoEXT extends VkGraphicsPipelineCreateInfo,VkComputePipelineCreateInfo,VkPipelineShaderStageCreateInfo,VkRayTracingPipelineCreateInfoKHR
pub struct PipelineRobustnessCreateInfoEXT {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    storage_buffers                              PipelineRobustnessBufferBehaviorEXT
    uniform_buffers                              PipelineRobustnessBufferBehaviorEXT
    vertex_inputs                                PipelineRobustnessBufferBehaviorEXT
    images                                       PipelineRobustnessImageBehaviorEXT
} 



// VK_EXT_conditional_rendering is a preprocessor guard. Do not pass it to API calls.
const ext_conditional_rendering = 1
pub const ext_conditional_rendering_spec_version = 2
pub const ext_conditional_rendering_extension_name = "VK_EXT_conditional_rendering"

pub enum ConditionalRenderingFlagBitsEXT {
    conditional_rendering_inverted_bit_ext = int(0x00000001)
    conditional_rendering_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type ConditionalRenderingFlagsEXT = u32
pub struct ConditionalRenderingBeginInfoEXT {
mut:
    s_type                                StructureType
    p_next                                voidptr
    buffer                                C.Buffer
    offset                                DeviceSize
    flags                                 ConditionalRenderingFlagsEXT
} 

// PhysicalDeviceConditionalRenderingFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceConditionalRenderingFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    conditional_rendering  Bool32
    inherited_conditional_rendering Bool32
} 

// CommandBufferInheritanceConditionalRenderingInfoEXT extends VkCommandBufferInheritanceInfo
pub struct CommandBufferInheritanceConditionalRenderingInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    conditional_rendering_enable Bool32
} 

type VkCmdBeginConditionalRenderingEXT = fn (     C.CommandBuffer,     &ConditionalRenderingBeginInfoEXT) 

pub fn cmd_begin_conditional_rendering_ext(
    command_buffer                                  C.CommandBuffer,
    p_conditional_rendering_begin                   &ConditionalRenderingBeginInfoEXT)  {
      f := VkCmdBeginConditionalRenderingEXT((*loader_p).get_sym('vkCmdBeginConditionalRenderingEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBeginConditionalRenderingEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    p_conditional_rendering_begin)
}


type VkCmdEndConditionalRenderingEXT = fn (     C.CommandBuffer) 

pub fn cmd_end_conditional_rendering_ext(
    command_buffer                                  C.CommandBuffer)  {
      f := VkCmdEndConditionalRenderingEXT((*loader_p).get_sym('vkCmdEndConditionalRenderingEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEndConditionalRenderingEXT': ${err}")
        return 
    })
    f(
    command_buffer)
}




// VK_NV_clip_space_w_scaling is a preprocessor guard. Do not pass it to API calls.
const nv_clip_space_w_scaling = 1
pub const nv_clip_space_w_scaling_spec_version = 1
pub const nv_clip_space_w_scaling_extension_name = "VK_NV_clip_space_w_scaling"
pub struct ViewportWScalingNV {
mut:
    xcoeff       f32
    ycoeff       f32
} 

// PipelineViewportWScalingStateCreateInfoNV extends VkPipelineViewportStateCreateInfo
pub struct PipelineViewportWScalingStateCreateInfoNV {
mut:
    s_type                             StructureType
    p_next                             voidptr
    viewport_w_scaling_enable          Bool32
    viewport_count                     u32
    p_viewport_w_scalings              &ViewportWScalingNV
} 

type VkCmdSetViewportWScalingNV = fn (     C.CommandBuffer,     u32,     u32,     &ViewportWScalingNV) 

pub fn cmd_set_viewport_w_scaling_nv(
    command_buffer                                  C.CommandBuffer,
    first_viewport                                  u32,
    viewport_count                                  u32,
    p_viewport_w_scalings                           &ViewportWScalingNV)  {
      f := VkCmdSetViewportWScalingNV((*loader_p).get_sym('vkCmdSetViewportWScalingNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetViewportWScalingNV': ${err}")
        return 
    })
    f(
    command_buffer,
    first_viewport,
    viewport_count,
    p_viewport_w_scalings)
}




// VK_EXT_direct_mode_display is a preprocessor guard. Do not pass it to API calls.
const ext_direct_mode_display = 1
pub const ext_direct_mode_display_spec_version = 1
pub const ext_direct_mode_display_extension_name = "VK_EXT_direct_mode_display"
type VkReleaseDisplayEXT = fn (     C.PhysicalDevice,     C.DisplayKHR) Result

pub fn release_display_ext(
    physical_device                                 C.PhysicalDevice,
    display                                         C.DisplayKHR) Result {
      f := VkReleaseDisplayEXT((*loader_p).get_sym('vkReleaseDisplayEXT'
    ) or { 
        println("Couldn't load symbol for 'vkReleaseDisplayEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    display)
}




// VK_EXT_acquire_xlib_display is a preprocessor guard. Do not pass it to API calls.
const ext_acquire_xlib_display = 1
pub const ext_acquire_xlib_display_spec_version = 1
pub const ext_acquire_xlib_display_extension_name = "VK_EXT_acquire_xlib_display"
type VkAcquireXlibDisplayEXT = fn (     C.PhysicalDevice,     &C.DisplayKHR,     C.DisplayKHR) Result

pub fn acquire_xlib_display_ext(
    physical_device                                 C.PhysicalDevice,
    dpy                                             &C.DisplayKHR,
    display                                         C.DisplayKHR) Result {
      f := VkAcquireXlibDisplayEXT((*loader_p).get_sym('vkAcquireXlibDisplayEXT'
    ) or { 
        println("Couldn't load symbol for 'vkAcquireXlibDisplayEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    dpy,
    display)
}


type VkGetRandROutputDisplayEXT = fn (     C.PhysicalDevice,     &C.DisplayKHR,     u32,     &C.DisplayKHR) Result

pub fn get_rand_r_output_display_ext(
    physical_device                                 C.PhysicalDevice,
    dpy                                             &C.DisplayKHR,
    rr_output                                       u32,
    p_display                                       &C.DisplayKHR) Result {
      f := VkGetRandROutputDisplayEXT((*loader_p).get_sym('vkGetRandROutputDisplayEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetRandROutputDisplayEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    dpy,
    rr_output,
    p_display)
}




// VK_EXT_display_surface_counter is a preprocessor guard. Do not pass it to API calls.
const ext_display_surface_counter = 1
pub const ext_display_surface_counter_spec_version = 1
pub const ext_display_surface_counter_extension_name = "VK_EXT_display_surface_counter"

pub enum SurfaceCounterFlagBitsEXT {
    surface_counter_vblank_bit_ext = int(0x00000001)
    surface_counter_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type SurfaceCounterFlagsEXT = u32
pub struct SurfaceCapabilities2EXT {
mut:
    s_type                               StructureType
    p_next                               voidptr
    min_image_count                      u32
    max_image_count                      u32
    current_extent                       Extent2D
    min_image_extent                     Extent2D
    max_image_extent                     Extent2D
    max_image_array_layers               u32
    supported_transforms                 SurfaceTransformFlagsKHR
    current_transform                    SurfaceTransformFlagBitsKHR
    supported_composite_alpha            CompositeAlphaFlagsKHR
    supported_usage_flags                ImageUsageFlags
    supported_surface_counters           SurfaceCounterFlagsEXT
} 

type VkGetPhysicalDeviceSurfaceCapabilities2EXT = fn (     C.PhysicalDevice,     C.SurfaceKHR,     &SurfaceCapabilities2EXT) Result

pub fn get_physical_device_surface_capabilities2_ext(
    physical_device                                 C.PhysicalDevice,
    surface                                         C.SurfaceKHR,
    p_surface_capabilities                          &SurfaceCapabilities2EXT) Result {
      f := VkGetPhysicalDeviceSurfaceCapabilities2EXT((*loader_p).get_sym('vkGetPhysicalDeviceSurfaceCapabilities2EXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSurfaceCapabilities2EXT': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    surface,
    p_surface_capabilities)
}




// VK_EXT_display_control is a preprocessor guard. Do not pass it to API calls.
const ext_display_control = 1
pub const ext_display_control_spec_version  = 1
pub const ext_display_control_extension_name = "VK_EXT_display_control"

pub enum DisplayPowerStateEXT {
    display_power_state_off_ext = int(0)
    display_power_state_suspend_ext = int(1)
    display_power_state_on_ext = int(2)
    display_power_state_max_enum_ext = int(0x7FFFFFFF)
}


pub enum DeviceEventTypeEXT {
    device_event_type_display_hotplug_ext = int(0)
    device_event_type_max_enum_ext = int(0x7FFFFFFF)
}


pub enum DisplayEventTypeEXT {
    display_event_type_first_pixel_out_ext = int(0)
    display_event_type_max_enum_ext = int(0x7FFFFFFF)
}

pub struct DisplayPowerInfoEXT {
mut:
    s_type                        StructureType
    p_next                        voidptr
    power_state                   DisplayPowerStateEXT
} 

pub struct DeviceEventInfoEXT {
mut:
    s_type                      StructureType
    p_next                      voidptr
    device_event                DeviceEventTypeEXT
} 

pub struct DisplayEventInfoEXT {
mut:
    s_type                       StructureType
    p_next                       voidptr
    display_event                DisplayEventTypeEXT
} 

// SwapchainCounterCreateInfoEXT extends VkSwapchainCreateInfoKHR
pub struct SwapchainCounterCreateInfoEXT {
mut:
    s_type                          StructureType
    p_next                          voidptr
    surface_counters                SurfaceCounterFlagsEXT
} 

type VkDisplayPowerControlEXT = fn (     C.Device,     C.DisplayKHR,     &DisplayPowerInfoEXT) Result

pub fn display_power_control_ext(
    device                                          C.Device,
    display                                         C.DisplayKHR,
    p_display_power_info                            &DisplayPowerInfoEXT) Result {
      f := VkDisplayPowerControlEXT((*loader_p).get_sym('vkDisplayPowerControlEXT'
    ) or { 
        println("Couldn't load symbol for 'vkDisplayPowerControlEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    display,
    p_display_power_info)
}


type VkRegisterDeviceEventEXT = fn (     C.Device,     &DeviceEventInfoEXT,     &AllocationCallbacks,     &C.Fence) Result

pub fn register_device_event_ext(
    device                                          C.Device,
    p_device_event_info                             &DeviceEventInfoEXT,
    p_allocator                                     &AllocationCallbacks,
    p_fence                                         &C.Fence) Result {
      f := VkRegisterDeviceEventEXT((*loader_p).get_sym('vkRegisterDeviceEventEXT'
    ) or { 
        println("Couldn't load symbol for 'vkRegisterDeviceEventEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_device_event_info,
    p_allocator,
    p_fence)
}


type VkRegisterDisplayEventEXT = fn (     C.Device,     C.DisplayKHR,     &DisplayEventInfoEXT,     &AllocationCallbacks,     &C.Fence) Result

pub fn register_display_event_ext(
    device                                          C.Device,
    display                                         C.DisplayKHR,
    p_display_event_info                            &DisplayEventInfoEXT,
    p_allocator                                     &AllocationCallbacks,
    p_fence                                         &C.Fence) Result {
      f := VkRegisterDisplayEventEXT((*loader_p).get_sym('vkRegisterDisplayEventEXT'
    ) or { 
        println("Couldn't load symbol for 'vkRegisterDisplayEventEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    display,
    p_display_event_info,
    p_allocator,
    p_fence)
}


type VkGetSwapchainCounterEXT = fn (     C.Device,     C.SwapchainKHR,     SurfaceCounterFlagBitsEXT,     &u64) Result

pub fn get_swapchain_counter_ext(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR,
    counter                                         SurfaceCounterFlagBitsEXT,
    p_counter_value                                 &u64) Result {
      f := VkGetSwapchainCounterEXT((*loader_p).get_sym('vkGetSwapchainCounterEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetSwapchainCounterEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain,
    counter,
    p_counter_value)
}




// VK_GOOGLE_display_timing is a preprocessor guard. Do not pass it to API calls.
const google_display_timing = 1
pub const google_display_timing_spec_version = 1
pub const google_display_timing_extension_name = "VK_GOOGE_display_timing"
pub struct RefreshCycleDurationGOOGLE {
mut:
    refresh_duration u64
} 

pub struct PastPresentationTimingGOOGLE {
mut:
    present_id      u32
    desired_present_time u64
    actual_present_time u64
    earliest_present_time u64
    present_margin  u64
} 

pub struct PresentTimeGOOGLE {
mut:
    present_id      u32
    desired_present_time u64
} 

// PresentTimesInfoGOOGLE extends VkPresentInfoKHR
pub struct PresentTimesInfoGOOGLE {
mut:
    s_type                            StructureType
    p_next                            voidptr
    swapchain_count                   u32
    p_times                           &PresentTimeGOOGLE
} 

type VkGetRefreshCycleDurationGOOGLE = fn (     C.Device,     C.SwapchainKHR,     &RefreshCycleDurationGOOGLE) Result

pub fn get_refresh_cycle_duration_google(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR,
    p_display_timing_properties                     &RefreshCycleDurationGOOGLE) Result {
      f := VkGetRefreshCycleDurationGOOGLE((*loader_p).get_sym('vkGetRefreshCycleDurationGOOGLE'
    ) or { 
        println("Couldn't load symbol for 'vkGetRefreshCycleDurationGOOGLE': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain,
    p_display_timing_properties)
}


type VkGetPastPresentationTimingGOOGLE = fn (     C.Device,     C.SwapchainKHR,     &u32,     &PastPresentationTimingGOOGLE) Result

pub fn get_past_presentation_timing_google(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR,
    p_presentation_timing_count                     &u32,
    p_presentation_timings                          &PastPresentationTimingGOOGLE) Result {
      f := VkGetPastPresentationTimingGOOGLE((*loader_p).get_sym('vkGetPastPresentationTimingGOOGLE'
    ) or { 
        println("Couldn't load symbol for 'vkGetPastPresentationTimingGOOGLE': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain,
    p_presentation_timing_count,
    p_presentation_timings)
}




// VK_NV_sample_mask_override_coverage is a preprocessor guard. Do not pass it to API calls.
const nv_sample_mask_override_coverage = 1
pub const nv_sample_mask_override_coverage_spec_version = 1
pub const nv_sample_mask_override_coverage_extension_name = "VK_NV_sample_mask_override_coverage"


// VK_NV_geometry_shader_passthrough is a preprocessor guard. Do not pass it to API calls.
const nv_geometry_shader_passthrough = 1
pub const nv_geometry_shader_passthrough_spec_version = 1
pub const nv_geometry_shader_passthrough_extension_name = "VK_NV_geometry_shader_passthrough"


// VK_NV_viewport_array2 is a preprocessor guard. Do not pass it to API calls.
const nv_viewport_array2 = 1
pub const nv_viewport_array_2_spec_version  = 1
pub const nv_viewport_array_2_extension_name = "VK_NV_viewport_array2"
pub const nv_viewport_array2_spec_version   = nv_viewport_array_2_spec_version
pub const nv_viewport_array2_extension_name = nv_viewport_array_2_extension_name


// VK_NVX_multiview_per_view_attributes is a preprocessor guard. Do not pass it to API calls.
const nvx_multiview_per_view_attributes = 1
pub const nvx_multiview_per_view_attributes_spec_version = 1
pub const nvx_multiview_per_view_attributes_extension_name = "VK_NVX_multiview_per_view_attributes"
// PhysicalDeviceMultiviewPerViewAttributesPropertiesNVX extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceMultiviewPerViewAttributesPropertiesNVX {
mut:
    s_type                 StructureType
    p_next                 voidptr
    per_view_position_all_components Bool32
} 



// VK_NV_viewport_swizzle is a preprocessor guard. Do not pass it to API calls.
const nv_viewport_swizzle = 1
pub const nv_viewport_swizzle_spec_version  = 1
pub const nv_viewport_swizzle_extension_name = "VK_NV_viewport_swizzle"

pub enum ViewportCoordinateSwizzleNV {
    viewport_coordinate_swizzle_positive_x_nv = int(0)
    viewport_coordinate_swizzle_negative_x_nv = int(1)
    viewport_coordinate_swizzle_positive_y_nv = int(2)
    viewport_coordinate_swizzle_negative_y_nv = int(3)
    viewport_coordinate_swizzle_positive_z_nv = int(4)
    viewport_coordinate_swizzle_negative_z_nv = int(5)
    viewport_coordinate_swizzle_positive_w_nv = int(6)
    viewport_coordinate_swizzle_negative_w_nv = int(7)
    viewport_coordinate_swizzle_max_enum_nv = int(0x7FFFFFFF)
}

pub type PipelineViewportSwizzleStateCreateFlagsNV = u32
pub struct ViewportSwizzleNV {
mut:
    x                                    ViewportCoordinateSwizzleNV
    y                                    ViewportCoordinateSwizzleNV
    z                                    ViewportCoordinateSwizzleNV
    w                                    ViewportCoordinateSwizzleNV
} 

// PipelineViewportSwizzleStateCreateInfoNV extends VkPipelineViewportStateCreateInfo
pub struct PipelineViewportSwizzleStateCreateInfoNV {
mut:
    s_type                                             StructureType
    p_next                                             voidptr
    flags                                              PipelineViewportSwizzleStateCreateFlagsNV
    viewport_count                                     u32
    p_viewport_swizzles                                &ViewportSwizzleNV
} 



// VK_EXT_discard_rectangles is a preprocessor guard. Do not pass it to API calls.
const ext_discard_rectangles = 1
pub const ext_discard_rectangles_spec_version = 2
pub const ext_discard_rectangles_extension_name = "VK_EXT_discard_rectangles"

pub enum DiscardRectangleModeEXT {
    discard_rectangle_mode_inclusive_ext = int(0)
    discard_rectangle_mode_exclusive_ext = int(1)
    discard_rectangle_mode_max_enum_ext = int(0x7FFFFFFF)
}

pub type PipelineDiscardRectangleStateCreateFlagsEXT = u32
// PhysicalDeviceDiscardRectanglePropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceDiscardRectanglePropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_discard_rectangles u32
} 

// PipelineDiscardRectangleStateCreateInfoEXT extends VkGraphicsPipelineCreateInfo
pub struct PipelineDiscardRectangleStateCreateInfoEXT {
mut:
    s_type                                               StructureType
    p_next                                               voidptr
    flags                                                PipelineDiscardRectangleStateCreateFlagsEXT
    discard_rectangle_mode                               DiscardRectangleModeEXT
    discard_rectangle_count                              u32
    p_discard_rectangles                                 &Rect2D
} 

type VkCmdSetDiscardRectangleEXT = fn (     C.CommandBuffer,     u32,     u32,     &Rect2D) 

pub fn cmd_set_discard_rectangle_ext(
    command_buffer                                  C.CommandBuffer,
    first_discard_rectangle                         u32,
    discard_rectangle_count                         u32,
    p_discard_rectangles                            &Rect2D)  {
      f := VkCmdSetDiscardRectangleEXT((*loader_p).get_sym('vkCmdSetDiscardRectangleEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDiscardRectangleEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    first_discard_rectangle,
    discard_rectangle_count,
    p_discard_rectangles)
}


type VkCmdSetDiscardRectangleEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_discard_rectangle_enable_ext(
    command_buffer                                  C.CommandBuffer,
    discard_rectangle_enable                        Bool32)  {
      f := VkCmdSetDiscardRectangleEnableEXT((*loader_p).get_sym('vkCmdSetDiscardRectangleEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDiscardRectangleEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    discard_rectangle_enable)
}


type VkCmdSetDiscardRectangleModeEXT = fn (     C.CommandBuffer,     DiscardRectangleModeEXT) 

pub fn cmd_set_discard_rectangle_mode_ext(
    command_buffer                                  C.CommandBuffer,
    discard_rectangle_mode                          DiscardRectangleModeEXT)  {
      f := VkCmdSetDiscardRectangleModeEXT((*loader_p).get_sym('vkCmdSetDiscardRectangleModeEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDiscardRectangleModeEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    discard_rectangle_mode)
}




// VK_EXT_conservative_rasterization is a preprocessor guard. Do not pass it to API calls.
const ext_conservative_rasterization = 1
pub const ext_conservative_rasterization_spec_version = 1
pub const ext_conservative_rasterization_extension_name = "VK_EXT_conservative_rasterization"

pub enum ConservativeRasterizationModeEXT {
    conservative_rasterization_mode_disabled_ext = int(0)
    conservative_rasterization_mode_overestimate_ext = int(1)
    conservative_rasterization_mode_underestimate_ext = int(2)
    conservative_rasterization_mode_max_enum_ext = int(0x7FFFFFFF)
}

pub type PipelineRasterizationConservativeStateCreateFlagsEXT = u32
// PhysicalDeviceConservativeRasterizationPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceConservativeRasterizationPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    primitive_overestimation_size f32
    max_extra_primitive_overestimation_size f32
    extra_primitive_overestimation_size_granularity f32
    primitive_underestimation Bool32
    conservative_point_and_line_rasterization Bool32
    degenerate_triangles_rasterized Bool32
    degenerate_lines_rasterized Bool32
    fully_covered_fragment_shader_input_variable Bool32
    conservative_rasterization_post_depth_coverage Bool32
} 

// PipelineRasterizationConservativeStateCreateInfoEXT extends VkPipelineRasterizationStateCreateInfo
pub struct PipelineRasterizationConservativeStateCreateInfoEXT {
mut:
    s_type                                                        StructureType
    p_next                                                        voidptr
    flags                                                         PipelineRasterizationConservativeStateCreateFlagsEXT
    conservative_rasterization_mode                               ConservativeRasterizationModeEXT
    extra_primitive_overestimation_size                           f32
} 



// VK_EXT_depth_clip_enable is a preprocessor guard. Do not pass it to API calls.
const ext_depth_clip_enable = 1
pub const ext_depth_clip_enable_spec_version = 1
pub const ext_depth_clip_enable_extension_name = "VK_EXT_depth_clip_enable"
pub type PipelineRasterizationDepthClipStateCreateFlagsEXT = u32
// PhysicalDeviceDepthClipEnableFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDepthClipEnableFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    depth_clip_enable      Bool32
} 

// PipelineRasterizationDepthClipStateCreateInfoEXT extends VkPipelineRasterizationStateCreateInfo
pub struct PipelineRasterizationDepthClipStateCreateInfoEXT {
mut:
    s_type                                                     StructureType
    p_next                                                     voidptr
    flags                                                      PipelineRasterizationDepthClipStateCreateFlagsEXT
    depth_clip_enable                                          Bool32
} 



// VK_EXT_swapchain_colorspace is a preprocessor guard. Do not pass it to API calls.
const ext_swapchain_colorspace = 1
pub const ext_swapchain_color_space_spec_version = 4
pub const ext_swapchain_color_space_extension_name = "VK_EXT_swapchain_colorspace"


// VK_EXT_hdr_metadata is a preprocessor guard. Do not pass it to API calls.
const ext_hdr_metadata = 1
pub const ext_hdr_metadata_spec_version     = 2
pub const ext_hdr_metadata_extension_name   = "VK_EXT_hdr_metadata"
pub struct XYColorEXT {
mut:
    x            f32
    y            f32
} 

pub struct HdrMetadataEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    display_primary_red    XYColorEXT
    display_primary_green  XYColorEXT
    display_primary_blue   XYColorEXT
    white_point            XYColorEXT
    max_luminance          f32
    min_luminance          f32
    max_content_light_level f32
    max_frame_average_light_level f32
} 

type VkSetHdrMetadataEXT = fn (     C.Device,     u32,     &C.SwapchainKHR,     &HdrMetadataEXT) 

pub fn set_hdr_metadata_ext(
    device                                          C.Device,
    swapchain_count                                 u32,
    p_swapchains                                    &C.SwapchainKHR,
    p_metadata                                      &HdrMetadataEXT)  {
      f := VkSetHdrMetadataEXT((*loader_p).get_sym('vkSetHdrMetadataEXT'
    ) or { 
        println("Couldn't load symbol for 'vkSetHdrMetadataEXT': ${err}")
        return 
    })
    f(
    device,
    swapchain_count,
    p_swapchains,
    p_metadata)
}




// VK_IMG_relaxed_line_rasterization is a preprocessor guard. Do not pass it to API calls.
const img_relaxed_line_rasterization = 1
pub const img_relaxed_line_rasterization_spec_version = 1
pub const img_relaxed_line_rasterization_extension_name = "VK_IMG_relaxed_line_rasterization"
// PhysicalDeviceRelaxedLineRasterizationFeaturesIMG extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRelaxedLineRasterizationFeaturesIMG {
mut:
    s_type                 StructureType
    p_next                 voidptr
    relaxed_line_rasterization Bool32
} 



// VK_MVK_ios_surface is a preprocessor guard. Do not pass it to API calls.
const mvk_ios_surface = 1
pub const mvk_ios_surface_spec_version      = 3
pub const mvk_ios_surface_extension_name    = "VK_MVK_ios_surface"
pub type IOSSurfaceCreateFlagsMVK = u32
pub struct IOSSurfaceCreateInfoMVK {
mut:
    s_type                            StructureType
    p_next                            voidptr
    flags                             IOSSurfaceCreateFlagsMVK
    p_view                            voidptr
} 

type VkCreateIOSSurfaceMVK = fn (     C.Instance,     &IOSSurfaceCreateInfoMVK,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_ios_surface_mvk(
    instance                                        C.Instance,
    p_create_info                                   &IOSSurfaceCreateInfoMVK,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateIOSSurfaceMVK((*loader_p).get_sym('vkCreateIOSSurfaceMVK'
    ) or { 
        println("Couldn't load symbol for 'vkCreateIOSSurfaceMVK': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}




// VK_MVK_macos_surface is a preprocessor guard. Do not pass it to API calls.
const mvk_macos_surface = 1
pub const mvk_macos_surface_spec_version    = 3
pub const mvk_macos_surface_extension_name  = "VK_MVK_macos_surface"
pub type MacOSSurfaceCreateFlagsMVK = u32
pub struct MacOSSurfaceCreateInfoMVK {
mut:
    s_type                              StructureType
    p_next                              voidptr
    flags                               MacOSSurfaceCreateFlagsMVK
    p_view                              voidptr
} 

type VkCreateMacOSSurfaceMVK = fn (     C.Instance,     &MacOSSurfaceCreateInfoMVK,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_mac_os_surface_mvk(
    instance                                        C.Instance,
    p_create_info                                   &MacOSSurfaceCreateInfoMVK,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateMacOSSurfaceMVK((*loader_p).get_sym('vkCreateMacOSSurfaceMVK'
    ) or { 
        println("Couldn't load symbol for 'vkCreateMacOSSurfaceMVK': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}




// VK_EXT_external_memory_dma_buf is a preprocessor guard. Do not pass it to API calls.
const ext_external_memory_dma_buf = 1
pub const ext_external_memory_dma_buf_spec_version = 1
pub const ext_external_memory_dma_buf_extension_name = "VK_EXT_external_memory_dma_buf"


// VK_EXT_queue_family_foreign is a preprocessor guard. Do not pass it to API calls.
const ext_queue_family_foreign = 1
pub const ext_queue_family_foreign_spec_version = 1
pub const ext_queue_family_foreign_extension_name = "VK_EXT_queue_family_foreign"
pub const queue_family_foreign_ext          = ~u32(2)


// VK_EXT_debug_utils is a preprocessor guard. Do not pass it to API calls.
const ext_debug_utils = 1
pub type C.DebugUtilsMessengerEXT = voidptr
pub const ext_debug_utils_spec_version      = 2
pub const ext_debug_utils_extension_name    = "VK_EXT_debug_utils"
pub type DebugUtilsMessengerCallbackDataFlagsEXT = u32

pub enum DebugUtilsMessageSeverityFlagBitsEXT {
    debug_utils_message_severity_verbose_bit_ext = int(0x00000001)
    debug_utils_message_severity_info_bit_ext = int(0x00000010)
    debug_utils_message_severity_warning_bit_ext = int(0x00000100)
    debug_utils_message_severity_error_bit_ext = int(0x00001000)
    debug_utils_message_severity_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}


pub enum DebugUtilsMessageTypeFlagBitsEXT {
    debug_utils_message_type_general_bit_ext = int(0x00000001)
    debug_utils_message_type_validation_bit_ext = int(0x00000002)
    debug_utils_message_type_performance_bit_ext = int(0x00000004)
    debug_utils_message_type_device_address_binding_bit_ext = int(0x00000008)
    debug_utils_message_type_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type DebugUtilsMessageTypeFlagsEXT = u32
pub type DebugUtilsMessageSeverityFlagsEXT = u32
pub type DebugUtilsMessengerCreateFlagsEXT = u32
pub struct DebugUtilsLabelEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    p_label_name           &char
    color                  []f32
} 

// DebugUtilsObjectNameInfoEXT extends VkPipelineShaderStageCreateInfo
pub struct DebugUtilsObjectNameInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    object_type            ObjectType
    object_handle          u64
    p_object_name          &char
} 

pub struct DebugUtilsMessengerCallbackDataEXT {
mut:
    s_type                                           StructureType
    p_next                                           voidptr
    flags                                            DebugUtilsMessengerCallbackDataFlagsEXT
    p_message_id_name                                &char
    message_id_number                                i32
    p_message                                        &char
    queue_label_count                                u32
    p_queue_labels                                   &DebugUtilsLabelEXT
    cmd_buf_label_count                              u32
    p_cmd_buf_labels                                 &DebugUtilsLabelEXT
    object_count                                     u32
    p_objects                                        &DebugUtilsObjectNameInfoEXT
} 

pub type PFN_vkDebugUtilsMessengerCallbackEXT = fn (   messageSeverity                   DebugUtilsMessageSeverityFlagBitsEXT,   messageTypes                      DebugUtilsMessageTypeFlagsEXT,   pCallbackData                     &DebugUtilsMessengerCallbackDataEXT,   pUserData                         voidptr) voidptr
// DebugUtilsMessengerCreateInfoEXT extends VkInstanceCreateInfo
pub struct DebugUtilsMessengerCreateInfoEXT {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    flags                                       DebugUtilsMessengerCreateFlagsEXT
    message_severity                            DebugUtilsMessageSeverityFlagsEXT
    message_type                                DebugUtilsMessageTypeFlagsEXT
    pfn_user_callback                           PFN_vkDebugUtilsMessengerCallbackEXT = unsafe { nil }
    p_user_data                                 voidptr
} 

pub struct DebugUtilsObjectTagInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    object_type            ObjectType
    object_handle          u64
    tag_name               u64
    tag_size               usize
    p_tag                  voidptr
} 

type VkSetDebugUtilsObjectNameEXT = fn (     C.Device,     &DebugUtilsObjectNameInfoEXT) Result

pub fn set_debug_utils_object_name_ext(
    device                                          C.Device,
    p_name_info                                     &DebugUtilsObjectNameInfoEXT) Result {
      f := VkSetDebugUtilsObjectNameEXT((*loader_p).get_sym('vkSetDebugUtilsObjectNameEXT'
    ) or { 
        println("Couldn't load symbol for 'vkSetDebugUtilsObjectNameEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_name_info)
}


type VkSetDebugUtilsObjectTagEXT = fn (     C.Device,     &DebugUtilsObjectTagInfoEXT) Result

pub fn set_debug_utils_object_tag_ext(
    device                                          C.Device,
    p_tag_info                                      &DebugUtilsObjectTagInfoEXT) Result {
      f := VkSetDebugUtilsObjectTagEXT((*loader_p).get_sym('vkSetDebugUtilsObjectTagEXT'
    ) or { 
        println("Couldn't load symbol for 'vkSetDebugUtilsObjectTagEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_tag_info)
}


type VkQueueBeginDebugUtilsLabelEXT = fn (     C.Queue,     &DebugUtilsLabelEXT) 

pub fn queue_begin_debug_utils_label_ext(
    queue                                           C.Queue,
    p_label_info                                    &DebugUtilsLabelEXT)  {
      f := VkQueueBeginDebugUtilsLabelEXT((*loader_p).get_sym('vkQueueBeginDebugUtilsLabelEXT'
    ) or { 
        println("Couldn't load symbol for 'vkQueueBeginDebugUtilsLabelEXT': ${err}")
        return 
    })
    f(
    queue,
    p_label_info)
}


type VkQueueEndDebugUtilsLabelEXT = fn (     C.Queue) 

pub fn queue_end_debug_utils_label_ext(
    queue                                           C.Queue)  {
      f := VkQueueEndDebugUtilsLabelEXT((*loader_p).get_sym('vkQueueEndDebugUtilsLabelEXT'
    ) or { 
        println("Couldn't load symbol for 'vkQueueEndDebugUtilsLabelEXT': ${err}")
        return 
    })
    f(
    queue)
}


type VkQueueInsertDebugUtilsLabelEXT = fn (     C.Queue,     &DebugUtilsLabelEXT) 

pub fn queue_insert_debug_utils_label_ext(
    queue                                           C.Queue,
    p_label_info                                    &DebugUtilsLabelEXT)  {
      f := VkQueueInsertDebugUtilsLabelEXT((*loader_p).get_sym('vkQueueInsertDebugUtilsLabelEXT'
    ) or { 
        println("Couldn't load symbol for 'vkQueueInsertDebugUtilsLabelEXT': ${err}")
        return 
    })
    f(
    queue,
    p_label_info)
}


type VkCmdBeginDebugUtilsLabelEXT = fn (     C.CommandBuffer,     &DebugUtilsLabelEXT) 

pub fn cmd_begin_debug_utils_label_ext(
    command_buffer                                  C.CommandBuffer,
    p_label_info                                    &DebugUtilsLabelEXT)  {
      f := VkCmdBeginDebugUtilsLabelEXT((*loader_p).get_sym('vkCmdBeginDebugUtilsLabelEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBeginDebugUtilsLabelEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    p_label_info)
}


type VkCmdEndDebugUtilsLabelEXT = fn (     C.CommandBuffer) 

pub fn cmd_end_debug_utils_label_ext(
    command_buffer                                  C.CommandBuffer)  {
      f := VkCmdEndDebugUtilsLabelEXT((*loader_p).get_sym('vkCmdEndDebugUtilsLabelEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdEndDebugUtilsLabelEXT': ${err}")
        return 
    })
    f(
    command_buffer)
}


type VkCmdInsertDebugUtilsLabelEXT = fn (     C.CommandBuffer,     &DebugUtilsLabelEXT) 

pub fn cmd_insert_debug_utils_label_ext(
    command_buffer                                  C.CommandBuffer,
    p_label_info                                    &DebugUtilsLabelEXT)  {
      f := VkCmdInsertDebugUtilsLabelEXT((*loader_p).get_sym('vkCmdInsertDebugUtilsLabelEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdInsertDebugUtilsLabelEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    p_label_info)
}


type VkCreateDebugUtilsMessengerEXT = fn (     C.Instance,     &DebugUtilsMessengerCreateInfoEXT,     &AllocationCallbacks,     &C.DebugUtilsMessengerEXT) Result

pub fn create_debug_utils_messenger_ext(
    instance                                        C.Instance,
    p_create_info                                   &DebugUtilsMessengerCreateInfoEXT,
    p_allocator                                     &AllocationCallbacks,
    p_messenger                                     &C.DebugUtilsMessengerEXT) Result {
      f := VkCreateDebugUtilsMessengerEXT((*loader_p).get_sym('vkCreateDebugUtilsMessengerEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCreateDebugUtilsMessengerEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_messenger)
}


type VkDestroyDebugUtilsMessengerEXT = fn (     C.Instance,     C.DebugUtilsMessengerEXT,     &AllocationCallbacks) 

pub fn destroy_debug_utils_messenger_ext(
    instance                                        C.Instance,
    messenger                                       C.DebugUtilsMessengerEXT,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyDebugUtilsMessengerEXT((*loader_p).get_sym('vkDestroyDebugUtilsMessengerEXT'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyDebugUtilsMessengerEXT': ${err}")
        return 
    })
    f(
    instance,
    messenger,
    p_allocator)
}


type VkSubmitDebugUtilsMessageEXT = fn (     C.Instance,     DebugUtilsMessageSeverityFlagBitsEXT,     DebugUtilsMessageTypeFlagsEXT,     &DebugUtilsMessengerCallbackDataEXT) 

pub fn submit_debug_utils_message_ext(
    instance                                        C.Instance,
    message_severity                                DebugUtilsMessageSeverityFlagBitsEXT,
    message_types                                   DebugUtilsMessageTypeFlagsEXT,
    p_callback_data                                 &DebugUtilsMessengerCallbackDataEXT)  {
      f := VkSubmitDebugUtilsMessageEXT((*loader_p).get_sym('vkSubmitDebugUtilsMessageEXT'
    ) or { 
        println("Couldn't load symbol for 'vkSubmitDebugUtilsMessageEXT': ${err}")
        return 
    })
    f(
    instance,
    message_severity,
    message_types,
    p_callback_data)
}




// VK_ANDROID_external_memory_android_hardware_buffer is a preprocessor guard. Do not pass it to API calls.
const android_external_memory_android_hardware_buffer = 1
pub const android_external_memory_android_hardware_buffer_spec_version = 5
pub const android_external_memory_android_hardware_buffer_extension_name = "VK_ANDROID_external_memory_android_hardware_buffer"
// AndroidHardwareBufferUsageANDROID extends VkImageFormatProperties2
pub struct AndroidHardwareBufferUsageANDROID {
mut:
    s_type                 StructureType
    p_next                 voidptr
    android_hardware_buffer_usage u64
} 

pub struct AndroidHardwareBufferPropertiesANDROID {
mut:
    s_type                 StructureType
    p_next                 voidptr
    allocation_size        DeviceSize
    memory_type_bits       u32
} 

// AndroidHardwareBufferFormatPropertiesANDROID extends VkAndroidHardwareBufferPropertiesANDROID
pub struct AndroidHardwareBufferFormatPropertiesANDROID {
mut:
    s_type                               StructureType
    p_next                               voidptr
    format                               Format
    external_format                      u64
    format_features                      FormatFeatureFlags
    sampler_ycbcr_conversion_components  ComponentMapping
    suggested_ycbcr_model                SamplerYcbcrModelConversion
    suggested_ycbcr_range                SamplerYcbcrRange
    suggested_x_chroma_offset            ChromaLocation
    suggested_y_chroma_offset            ChromaLocation
} 

// ImportAndroidHardwareBufferInfoANDROID extends VkMemoryAllocateInfo
pub struct ImportAndroidHardwareBufferInfoANDROID {
mut:
    s_type                         StructureType
    p_next                         voidptr
    buffer                         voidptr
} 

pub struct MemoryGetAndroidHardwareBufferInfoANDROID {
mut:
    s_type                 StructureType
    p_next                 voidptr
    memory                 C.DeviceMemory
} 

// ExternalFormatANDROID extends VkImageCreateInfo,VkSamplerYcbcrConversionCreateInfo,VkAttachmentDescription2,VkGraphicsPipelineCreateInfo,VkCommandBufferInheritanceInfo
pub struct ExternalFormatANDROID {
mut:
    s_type                 StructureType
    p_next                 voidptr
    external_format        u64
} 

// AndroidHardwareBufferFormatProperties2ANDROID extends VkAndroidHardwareBufferPropertiesANDROID
pub struct AndroidHardwareBufferFormatProperties2ANDROID {
mut:
    s_type                               StructureType
    p_next                               voidptr
    format                               Format
    external_format                      u64
    format_features                      FormatFeatureFlags2
    sampler_ycbcr_conversion_components  ComponentMapping
    suggested_ycbcr_model                SamplerYcbcrModelConversion
    suggested_ycbcr_range                SamplerYcbcrRange
    suggested_x_chroma_offset            ChromaLocation
    suggested_y_chroma_offset            ChromaLocation
} 

type VkGetAndroidHardwareBufferPropertiesANDROID = fn (     C.Device,     voidptr,     &AndroidHardwareBufferPropertiesANDROID) Result

pub fn get_android_hardware_buffer_properties_android(
    device                                          C.Device,
    buffer                                          voidptr,
    p_properties                                    &AndroidHardwareBufferPropertiesANDROID) Result {
      f := VkGetAndroidHardwareBufferPropertiesANDROID((*loader_p).get_sym('vkGetAndroidHardwareBufferPropertiesANDROID'
    ) or { 
        println("Couldn't load symbol for 'vkGetAndroidHardwareBufferPropertiesANDROID': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    buffer,
    p_properties)
}


type VkGetMemoryAndroidHardwareBufferANDROID = fn (     C.Device,     &MemoryGetAndroidHardwareBufferInfoANDROID,     voidptr) Result

pub fn get_memory_android_hardware_buffer_android(
    device                                          C.Device,
    p_info                                          &MemoryGetAndroidHardwareBufferInfoANDROID,
    p_buffer                                        voidptr) Result {
      f := VkGetMemoryAndroidHardwareBufferANDROID((*loader_p).get_sym('vkGetMemoryAndroidHardwareBufferANDROID'
    ) or { 
        println("Couldn't load symbol for 'vkGetMemoryAndroidHardwareBufferANDROID': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_info,
    p_buffer)
}




// VK_EXT_sampler_filter_minmax is a preprocessor guard. Do not pass it to API calls.
const ext_sampler_filter_minmax = 1
pub const ext_sampler_filter_minmax_spec_version = 2
pub const ext_sampler_filter_minmax_extension_name = "VK_EXT_sampler_filter_minmax"
pub type SamplerReductionModeEXT = SamplerReductionMode

pub type SamplerReductionModeCreateInfoEXT = SamplerReductionModeCreateInfo

pub type PhysicalDeviceSamplerFilterMinmaxPropertiesEXT = PhysicalDeviceSamplerFilterMinmaxProperties



// VK_AMD_gpu_shader_int16 is a preprocessor guard. Do not pass it to API calls.
const amd_gpu_shader_int16 = 1
pub const amd_gpu_shader_int16_spec_version = 2
pub const amd_gpu_shader_int16_extension_name = "VK_AMD_gpu_shader_int16"


// VK_AMDX_shader_enqueue is a preprocessor guard. Do not pass it to API calls.
const amdx_shader_enqueue = 1
pub const amdx_shader_enqueue_spec_version  = 1
pub const amdx_shader_enqueue_extension_name = "VK_AMDX_shader_enqueue"
pub const shader_index_unused_amdx          = ~u32(0)
// PhysicalDeviceShaderEnqueueFeaturesAMDX extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderEnqueueFeaturesAMDX {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_enqueue         Bool32
} 

// PhysicalDeviceShaderEnqueuePropertiesAMDX extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceShaderEnqueuePropertiesAMDX {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_execution_graph_depth u32
    max_execution_graph_shader_output_nodes u32
    max_execution_graph_shader_payload_size u32
    max_execution_graph_shader_payload_count u32
    execution_graph_dispatch_address_alignment u32
} 

pub struct ExecutionGraphPipelineScratchSizeAMDX {
mut:
    s_type                 StructureType
    p_next                 voidptr
    size                   DeviceSize
} 

pub struct ExecutionGraphPipelineCreateInfoAMDX {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    flags                                         PipelineCreateFlags
    stage_count                                   u32
    p_stages                                      &PipelineShaderStageCreateInfo
    p_library_info                                &PipelineLibraryCreateInfoKHR
    layout                                        C.PipelineLayout
    base_pipeline_handle                          C.Pipeline
    base_pipeline_index                           i32
} 

pub union DeviceOrHostAddressConstAMDX {
mut:
    device_address         DeviceAddress
    host_address           voidptr
} 

pub struct DispatchGraphInfoAMDX {
mut:
    node_index                            u32
    payload_count                         u32
    payloads                              DeviceOrHostAddressConstAMDX
    payload_stride                        u64
} 

pub struct DispatchGraphCountInfoAMDX {
mut:
    count                                 u32
    infos                                 DeviceOrHostAddressConstAMDX
    stride                                u64
} 

// PipelineShaderStageNodeCreateInfoAMDX extends VkPipelineShaderStageCreateInfo
pub struct PipelineShaderStageNodeCreateInfoAMDX {
mut:
    s_type                   StructureType
    p_next                   voidptr
    p_name                   &char
    index                    u32
} 

type VkCreateExecutionGraphPipelinesAMDX = fn (     C.Device,     C.PipelineCache,     u32,     &ExecutionGraphPipelineCreateInfoAMDX,     &AllocationCallbacks,     &C.Pipeline) Result

pub fn create_execution_graph_pipelines_amdx(
    device                                          C.Device,
    pipeline_cache                                  C.PipelineCache,
    create_info_count                               u32,
    p_create_infos                                  &ExecutionGraphPipelineCreateInfoAMDX,
    p_allocator                                     &AllocationCallbacks,
    p_pipelines                                     &C.Pipeline) Result {
      f := VkCreateExecutionGraphPipelinesAMDX((*loader_p).get_sym('vkCreateExecutionGraphPipelinesAMDX'
    ) or { 
        println("Couldn't load symbol for 'vkCreateExecutionGraphPipelinesAMDX': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    pipeline_cache,
    create_info_count,
    p_create_infos,
    p_allocator,
    p_pipelines)
}


type VkGetExecutionGraphPipelineScratchSizeAMDX = fn (     C.Device,     C.Pipeline,     &ExecutionGraphPipelineScratchSizeAMDX) Result

pub fn get_execution_graph_pipeline_scratch_size_amdx(
    device                                          C.Device,
    execution_graph                                 C.Pipeline,
    p_size_info                                     &ExecutionGraphPipelineScratchSizeAMDX) Result {
      f := VkGetExecutionGraphPipelineScratchSizeAMDX((*loader_p).get_sym('vkGetExecutionGraphPipelineScratchSizeAMDX'
    ) or { 
        println("Couldn't load symbol for 'vkGetExecutionGraphPipelineScratchSizeAMDX': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    execution_graph,
    p_size_info)
}


type VkGetExecutionGraphPipelineNodeIndexAMDX = fn (     C.Device,     C.Pipeline,     &PipelineShaderStageNodeCreateInfoAMDX,     &u32) Result

pub fn get_execution_graph_pipeline_node_index_amdx(
    device                                          C.Device,
    execution_graph                                 C.Pipeline,
    p_node_info                                     &PipelineShaderStageNodeCreateInfoAMDX,
    p_node_index                                    &u32) Result {
      f := VkGetExecutionGraphPipelineNodeIndexAMDX((*loader_p).get_sym('vkGetExecutionGraphPipelineNodeIndexAMDX'
    ) or { 
        println("Couldn't load symbol for 'vkGetExecutionGraphPipelineNodeIndexAMDX': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    execution_graph,
    p_node_info,
    p_node_index)
}


type VkCmdInitializeGraphScratchMemoryAMDX = fn (     C.CommandBuffer,     DeviceAddress) 

pub fn cmd_initialize_graph_scratch_memory_amdx(
    command_buffer                                  C.CommandBuffer,
    scratch                                         DeviceAddress)  {
      f := VkCmdInitializeGraphScratchMemoryAMDX((*loader_p).get_sym('vkCmdInitializeGraphScratchMemoryAMDX'
    ) or { 
        println("Couldn't load symbol for 'vkCmdInitializeGraphScratchMemoryAMDX': ${err}")
        return 
    })
    f(
    command_buffer,
    scratch)
}


type VkCmdDispatchGraphAMDX = fn (     C.CommandBuffer,     DeviceAddress,     &DispatchGraphCountInfoAMDX) 

pub fn cmd_dispatch_graph_amdx(
    command_buffer                                  C.CommandBuffer,
    scratch                                         DeviceAddress,
    p_count_info                                    &DispatchGraphCountInfoAMDX)  {
      f := VkCmdDispatchGraphAMDX((*loader_p).get_sym('vkCmdDispatchGraphAMDX'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDispatchGraphAMDX': ${err}")
        return 
    })
    f(
    command_buffer,
    scratch,
    p_count_info)
}


type VkCmdDispatchGraphIndirectAMDX = fn (     C.CommandBuffer,     DeviceAddress,     &DispatchGraphCountInfoAMDX) 

pub fn cmd_dispatch_graph_indirect_amdx(
    command_buffer                                  C.CommandBuffer,
    scratch                                         DeviceAddress,
    p_count_info                                    &DispatchGraphCountInfoAMDX)  {
      f := VkCmdDispatchGraphIndirectAMDX((*loader_p).get_sym('vkCmdDispatchGraphIndirectAMDX'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDispatchGraphIndirectAMDX': ${err}")
        return 
    })
    f(
    command_buffer,
    scratch,
    p_count_info)
}


type VkCmdDispatchGraphIndirectCountAMDX = fn (     C.CommandBuffer,     DeviceAddress,     DeviceAddress) 

pub fn cmd_dispatch_graph_indirect_count_amdx(
    command_buffer                                  C.CommandBuffer,
    scratch                                         DeviceAddress,
    count_info                                      DeviceAddress)  {
      f := VkCmdDispatchGraphIndirectCountAMDX((*loader_p).get_sym('vkCmdDispatchGraphIndirectCountAMDX'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDispatchGraphIndirectCountAMDX': ${err}")
        return 
    })
    f(
    command_buffer,
    scratch,
    count_info)
}




// VK_AMD_mixed_attachment_samples is a preprocessor guard. Do not pass it to API calls.
const amd_mixed_attachment_samples = 1
pub const amd_mixed_attachment_samples_spec_version = 1
pub const amd_mixed_attachment_samples_extension_name = "VK_AMD_mixed_attachment_samples"


// VK_AMD_shader_fragment_mask is a preprocessor guard. Do not pass it to API calls.
const amd_shader_fragment_mask = 1
pub const amd_shader_fragment_mask_spec_version = 1
pub const amd_shader_fragment_mask_extension_name = "VK_AMD_shader_fragment_mask"


// VK_EXT_inline_uniform_block is a preprocessor guard. Do not pass it to API calls.
const ext_inline_uniform_block = 1
pub const ext_inline_uniform_block_spec_version = 1
pub const ext_inline_uniform_block_extension_name = "VK_EXT_inline_uniform_block"
pub type PhysicalDeviceInlineUniformBlockFeaturesEXT = PhysicalDeviceInlineUniformBlockFeatures

pub type PhysicalDeviceInlineUniformBlockPropertiesEXT = PhysicalDeviceInlineUniformBlockProperties

pub type WriteDescriptorSetInlineUniformBlockEXT = WriteDescriptorSetInlineUniformBlock

pub type DescriptorPoolInlineUniformBlockCreateInfoEXT = DescriptorPoolInlineUniformBlockCreateInfo



// VK_EXT_shader_stencil_export is a preprocessor guard. Do not pass it to API calls.
const ext_shader_stencil_export = 1
pub const ext_shader_stencil_export_spec_version = 1
pub const ext_shader_stencil_export_extension_name = "VK_EXT_shader_stencil_export"


// VK_EXT_sample_locations is a preprocessor guard. Do not pass it to API calls.
const ext_sample_locations = 1
pub const ext_sample_locations_spec_version = 1
pub const ext_sample_locations_extension_name = "VK_EXT_sample_locations"
pub struct SampleLocationEXT {
mut:
    x            f32
    y            f32
} 

// SampleLocationsInfoEXT extends VkImageMemoryBarrier,VkImageMemoryBarrier2
pub struct SampleLocationsInfoEXT {
mut:
    s_type                            StructureType
    p_next                            voidptr
    sample_locations_per_pixel        SampleCountFlagBits
    sample_location_grid_size         Extent2D
    sample_locations_count            u32
    p_sample_locations                &SampleLocationEXT
} 

pub struct AttachmentSampleLocationsEXT {
mut:
    attachment_index                u32
    sample_locations_info           SampleLocationsInfoEXT
} 

pub struct SubpassSampleLocationsEXT {
mut:
    subpass_index                   u32
    sample_locations_info           SampleLocationsInfoEXT
} 

// RenderPassSampleLocationsBeginInfoEXT extends VkRenderPassBeginInfo
pub struct RenderPassSampleLocationsBeginInfoEXT {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    attachment_initial_sample_locations_count    u32
    p_attachment_initial_sample_locations        &AttachmentSampleLocationsEXT
    post_subpass_sample_locations_count          u32
    p_post_subpass_sample_locations              &SubpassSampleLocationsEXT
} 

// PipelineSampleLocationsStateCreateInfoEXT extends VkPipelineMultisampleStateCreateInfo
pub struct PipelineSampleLocationsStateCreateInfoEXT {
mut:
    s_type                          StructureType
    p_next                          voidptr
    sample_locations_enable         Bool32
    sample_locations_info           SampleLocationsInfoEXT
} 

// PhysicalDeviceSampleLocationsPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceSampleLocationsPropertiesEXT {
mut:
    s_type                    StructureType
    p_next                    voidptr
    sample_location_sample_counts SampleCountFlags
    max_sample_location_grid_size Extent2D
    sample_location_coordinate_range []f32
    sample_location_sub_pixel_bits u32
    variable_sample_locations Bool32
} 

pub struct MultisamplePropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_sample_location_grid_size Extent2D
} 

type VkCmdSetSampleLocationsEXT = fn (     C.CommandBuffer,     &SampleLocationsInfoEXT) 

pub fn cmd_set_sample_locations_ext(
    command_buffer                                  C.CommandBuffer,
    p_sample_locations_info                         &SampleLocationsInfoEXT)  {
      f := VkCmdSetSampleLocationsEXT((*loader_p).get_sym('vkCmdSetSampleLocationsEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetSampleLocationsEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    p_sample_locations_info)
}


type VkGetPhysicalDeviceMultisamplePropertiesEXT = fn (     C.PhysicalDevice,     SampleCountFlagBits,     &MultisamplePropertiesEXT) 

pub fn get_physical_device_multisample_properties_ext(
    physical_device                                 C.PhysicalDevice,
    samples                                         SampleCountFlagBits,
    p_multisample_properties                        &MultisamplePropertiesEXT)  {
      f := VkGetPhysicalDeviceMultisamplePropertiesEXT((*loader_p).get_sym('vkGetPhysicalDeviceMultisamplePropertiesEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceMultisamplePropertiesEXT': ${err}")
        return 
    })
    f(
    physical_device,
    samples,
    p_multisample_properties)
}




// VK_EXT_blend_operation_advanced is a preprocessor guard. Do not pass it to API calls.
const ext_blend_operation_advanced = 1
pub const ext_blend_operation_advanced_spec_version = 2
pub const ext_blend_operation_advanced_extension_name = "VK_EXT_blend_operation_advanced"

pub enum BlendOverlapEXT {
    blend_overlap_uncorrelated_ext = int(0)
    blend_overlap_disjoint_ext = int(1)
    blend_overlap_conjoint_ext = int(2)
    blend_overlap_max_enum_ext = int(0x7FFFFFFF)
}

// PhysicalDeviceBlendOperationAdvancedFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceBlendOperationAdvancedFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    advanced_blend_coherent_operations Bool32
} 

// PhysicalDeviceBlendOperationAdvancedPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceBlendOperationAdvancedPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    advanced_blend_max_color_attachments u32
    advanced_blend_independent_blend Bool32
    advanced_blend_non_premultiplied_src_color Bool32
    advanced_blend_non_premultiplied_dst_color Bool32
    advanced_blend_correlated_overlap Bool32
    advanced_blend_all_operations Bool32
} 

// PipelineColorBlendAdvancedStateCreateInfoEXT extends VkPipelineColorBlendStateCreateInfo
pub struct PipelineColorBlendAdvancedStateCreateInfoEXT {
mut:
    s_type                   StructureType
    p_next                   voidptr
    src_premultiplied        Bool32
    dst_premultiplied        Bool32
    blend_overlap            BlendOverlapEXT
} 



// VK_NV_fragment_coverage_to_color is a preprocessor guard. Do not pass it to API calls.
const nv_fragment_coverage_to_color = 1
pub const nv_fragment_coverage_to_color_spec_version = 1
pub const nv_fragment_coverage_to_color_extension_name = "VK_NV_fragment_coverage_to_color"
pub type PipelineCoverageToColorStateCreateFlagsNV = u32
// PipelineCoverageToColorStateCreateInfoNV extends VkPipelineMultisampleStateCreateInfo
pub struct PipelineCoverageToColorStateCreateInfoNV {
mut:
    s_type                                             StructureType
    p_next                                             voidptr
    flags                                              PipelineCoverageToColorStateCreateFlagsNV
    coverage_to_color_enable                           Bool32
    coverage_to_color_location                         u32
} 



// VK_NV_framebuffer_mixed_samples is a preprocessor guard. Do not pass it to API calls.
const nv_framebuffer_mixed_samples = 1
pub const nv_framebuffer_mixed_samples_spec_version = 1
pub const nv_framebuffer_mixed_samples_extension_name = "VK_NV_framebuffer_mixed_samples"

pub enum CoverageModulationModeNV {
    coverage_modulation_mode_none_nv = int(0)
    coverage_modulation_mode_rgb_nv = int(1)
    coverage_modulation_mode_alpha_nv = int(2)
    coverage_modulation_mode_rgba_nv = int(3)
    coverage_modulation_mode_max_enum_nv = int(0x7FFFFFFF)
}

pub type PipelineCoverageModulationStateCreateFlagsNV = u32
// PipelineCoverageModulationStateCreateInfoNV extends VkPipelineMultisampleStateCreateInfo
pub struct PipelineCoverageModulationStateCreateInfoNV {
mut:
    s_type                                                StructureType
    p_next                                                voidptr
    flags                                                 PipelineCoverageModulationStateCreateFlagsNV
    coverage_modulation_mode                              CoverageModulationModeNV
    coverage_modulation_table_enable                      Bool32
    coverage_modulation_table_count                       u32
    p_coverage_modulation_table                           &f32
} 



// VK_NV_fill_rectangle is a preprocessor guard. Do not pass it to API calls.
const nv_fill_rectangle = 1
pub const nv_fill_rectangle_spec_version    = 1
pub const nv_fill_rectangle_extension_name  = "VK_NV_fill_rectangle"


// VK_NV_shader_sm_builtins is a preprocessor guard. Do not pass it to API calls.
const nv_shader_sm_builtins = 1
pub const nv_shader_sm_builtins_spec_version = 1
pub const nv_shader_sm_builtins_extension_name = "VK_NV_shader_sm_builtins"
// PhysicalDeviceShaderSMBuiltinsPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceShaderSMBuiltinsPropertiesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_sm_count        u32
    shader_warps_per_sm    u32
} 

// PhysicalDeviceShaderSMBuiltinsFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderSMBuiltinsFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_sm_builtins     Bool32
} 



// VK_EXT_post_depth_coverage is a preprocessor guard. Do not pass it to API calls.
const ext_post_depth_coverage = 1
pub const ext_post_depth_coverage_spec_version = 1
pub const ext_post_depth_coverage_extension_name = "VK_EXT_post_depth_coverage"


// VK_EXT_image_drm_format_modifier is a preprocessor guard. Do not pass it to API calls.
const ext_image_drm_format_modifier = 1
pub const ext_image_drm_format_modifier_spec_version = 2
pub const ext_image_drm_format_modifier_extension_name = "VK_EXT_image_drm_format_modifier"
pub struct DrmFormatModifierPropertiesEXT {
mut:
    drm_format_modifier         u64
    drm_format_modifier_plane_count u32
    drm_format_modifier_tiling_features FormatFeatureFlags
} 

// DrmFormatModifierPropertiesListEXT extends VkFormatProperties2
pub struct DrmFormatModifierPropertiesListEXT {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    drm_format_modifier_count                u32
    p_drm_format_modifier_properties         &DrmFormatModifierPropertiesEXT
} 

// PhysicalDeviceImageDrmFormatModifierInfoEXT extends VkPhysicalDeviceImageFormatInfo2
pub struct PhysicalDeviceImageDrmFormatModifierInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    drm_format_modifier    u64
    sharing_mode           SharingMode
    queue_family_index_count u32
    p_queue_family_indices &u32
} 

// ImageDrmFormatModifierListCreateInfoEXT extends VkImageCreateInfo
pub struct ImageDrmFormatModifierListCreateInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    drm_format_modifier_count u32
    p_drm_format_modifiers &u64
} 

// ImageDrmFormatModifierExplicitCreateInfoEXT extends VkImageCreateInfo
pub struct ImageDrmFormatModifierExplicitCreateInfoEXT {
mut:
    s_type                            StructureType
    p_next                            voidptr
    drm_format_modifier               u64
    drm_format_modifier_plane_count   u32
    p_plane_layouts                   &SubresourceLayout
} 

pub struct ImageDrmFormatModifierPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    drm_format_modifier    u64
} 

pub struct DrmFormatModifierProperties2EXT {
mut:
    drm_format_modifier          u64
    drm_format_modifier_plane_count u32
    drm_format_modifier_tiling_features FormatFeatureFlags2
} 

// DrmFormatModifierPropertiesList2EXT extends VkFormatProperties2
pub struct DrmFormatModifierPropertiesList2EXT {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    drm_format_modifier_count                 u32
    p_drm_format_modifier_properties          &DrmFormatModifierProperties2EXT
} 

type VkGetImageDrmFormatModifierPropertiesEXT = fn (     C.Device,     C.Image,     &ImageDrmFormatModifierPropertiesEXT) Result

pub fn get_image_drm_format_modifier_properties_ext(
    device                                          C.Device,
    image                                           C.Image,
    p_properties                                    &ImageDrmFormatModifierPropertiesEXT) Result {
      f := VkGetImageDrmFormatModifierPropertiesEXT((*loader_p).get_sym('vkGetImageDrmFormatModifierPropertiesEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageDrmFormatModifierPropertiesEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    image,
    p_properties)
}




// VK_EXT_validation_cache is a preprocessor guard. Do not pass it to API calls.
const ext_validation_cache = 1
pub type C.ValidationCacheEXT = voidptr
pub const ext_validation_cache_spec_version = 1
pub const ext_validation_cache_extension_name = "VK_EXT_validation_cache"

pub enum ValidationCacheHeaderVersionEXT {
    validation_cache_header_version_one_ext = int(1)
    validation_cache_header_version_max_enum_ext = int(0x7FFFFFFF)
}

pub type ValidationCacheCreateFlagsEXT = u32
pub struct ValidationCacheCreateInfoEXT {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    flags                                  ValidationCacheCreateFlagsEXT
    initial_data_size                      usize
    p_initial_data                         voidptr
} 

// ShaderModuleValidationCacheCreateInfoEXT extends VkShaderModuleCreateInfo,VkPipelineShaderStageCreateInfo
pub struct ShaderModuleValidationCacheCreateInfoEXT {
mut:
    s_type                      StructureType
    p_next                      voidptr
    validation_cache            C.ValidationCacheEXT
} 

type VkCreateValidationCacheEXT = fn (     C.Device,     &ValidationCacheCreateInfoEXT,     &AllocationCallbacks,     &C.ValidationCacheEXT) Result

pub fn create_validation_cache_ext(
    device                                          C.Device,
    p_create_info                                   &ValidationCacheCreateInfoEXT,
    p_allocator                                     &AllocationCallbacks,
    p_validation_cache                              &C.ValidationCacheEXT) Result {
      f := VkCreateValidationCacheEXT((*loader_p).get_sym('vkCreateValidationCacheEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCreateValidationCacheEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_validation_cache)
}


type VkDestroyValidationCacheEXT = fn (     C.Device,     C.ValidationCacheEXT,     &AllocationCallbacks) 

pub fn destroy_validation_cache_ext(
    device                                          C.Device,
    validation_cache                                C.ValidationCacheEXT,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyValidationCacheEXT((*loader_p).get_sym('vkDestroyValidationCacheEXT'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyValidationCacheEXT': ${err}")
        return 
    })
    f(
    device,
    validation_cache,
    p_allocator)
}


type VkMergeValidationCachesEXT = fn (     C.Device,     C.ValidationCacheEXT,     u32,     &C.ValidationCacheEXT) Result

pub fn merge_validation_caches_ext(
    device                                          C.Device,
    dst_cache                                       C.ValidationCacheEXT,
    src_cache_count                                 u32,
    p_src_caches                                    &C.ValidationCacheEXT) Result {
      f := VkMergeValidationCachesEXT((*loader_p).get_sym('vkMergeValidationCachesEXT'
    ) or { 
        println("Couldn't load symbol for 'vkMergeValidationCachesEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    dst_cache,
    src_cache_count,
    p_src_caches)
}


type VkGetValidationCacheDataEXT = fn (     C.Device,     C.ValidationCacheEXT,     &usize,     voidptr) Result

pub fn get_validation_cache_data_ext(
    device                                          C.Device,
    validation_cache                                C.ValidationCacheEXT,
    p_data_size                                     &usize,
    p_data                                          voidptr) Result {
      f := VkGetValidationCacheDataEXT((*loader_p).get_sym('vkGetValidationCacheDataEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetValidationCacheDataEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    validation_cache,
    p_data_size,
    p_data)
}




// VK_EXT_descriptor_indexing is a preprocessor guard. Do not pass it to API calls.
const ext_descriptor_indexing = 1
pub const ext_descriptor_indexing_spec_version = 2
pub const ext_descriptor_indexing_extension_name = "VK_EXT_descriptor_indexing"
pub type DescriptorBindingFlagBitsEXT = DescriptorBindingFlagBits

pub type DescriptorSetLayoutBindingFlagsCreateInfoEXT = DescriptorSetLayoutBindingFlagsCreateInfo

pub type PhysicalDeviceDescriptorIndexingFeaturesEXT = PhysicalDeviceDescriptorIndexingFeatures

pub type PhysicalDeviceDescriptorIndexingPropertiesEXT = PhysicalDeviceDescriptorIndexingProperties

pub type DescriptorSetVariableDescriptorCountAllocateInfoEXT = DescriptorSetVariableDescriptorCountAllocateInfo

pub type DescriptorSetVariableDescriptorCountLayoutSupportEXT = DescriptorSetVariableDescriptorCountLayoutSupport



// VK_EXT_shader_viewport_index_layer is a preprocessor guard. Do not pass it to API calls.
const ext_shader_viewport_index_layer = 1
pub const ext_shader_viewport_index_layer_spec_version = 1
pub const ext_shader_viewport_index_layer_extension_name = "VK_EXT_shader_viewport_index_layer"


// VK_NV_shading_rate_image is a preprocessor guard. Do not pass it to API calls.
const nv_shading_rate_image = 1
pub const nv_shading_rate_image_spec_version = 3
pub const nv_shading_rate_image_extension_name = "VK_NV_shading_rate_image"

pub enum ShadingRatePaletteEntryNV {
    shading_rate_palette_entry_no_invocations_nv = int(0)
    shading_rate_palette_entry_16_invocations_per_pixel_nv = int(1)
    shading_rate_palette_entry_8_invocations_per_pixel_nv = int(2)
    shading_rate_palette_entry_4_invocations_per_pixel_nv = int(3)
    shading_rate_palette_entry_2_invocations_per_pixel_nv = int(4)
    shading_rate_palette_entry_1_invocation_per_pixel_nv = int(5)
    shading_rate_palette_entry_1_invocation_per_2x1_pixels_nv = int(6)
    shading_rate_palette_entry_1_invocation_per_1x2_pixels_nv = int(7)
    shading_rate_palette_entry_1_invocation_per_2x2_pixels_nv = int(8)
    shading_rate_palette_entry_1_invocation_per_4x2_pixels_nv = int(9)
    shading_rate_palette_entry_1_invocation_per_2x4_pixels_nv = int(10)
    shading_rate_palette_entry_1_invocation_per_4x4_pixels_nv = int(11)
    shading_rate_palette_entry_max_enum_nv = int(0x7FFFFFFF)
}


pub enum CoarseSampleOrderTypeNV {
    coarse_sample_order_type_default_nv = int(0)
    coarse_sample_order_type_custom_nv = int(1)
    coarse_sample_order_type_pixel_major_nv = int(2)
    coarse_sample_order_type_sample_major_nv = int(3)
    coarse_sample_order_type_max_enum_nv = int(0x7FFFFFFF)
}

pub struct ShadingRatePaletteNV {
mut:
    shading_rate_palette_entry_count          u32
    p_shading_rate_palette_entries            &ShadingRatePaletteEntryNV
} 

// PipelineViewportShadingRateImageStateCreateInfoNV extends VkPipelineViewportStateCreateInfo
pub struct PipelineViewportShadingRateImageStateCreateInfoNV {
mut:
    s_type                               StructureType
    p_next                               voidptr
    shading_rate_image_enable            Bool32
    viewport_count                       u32
    p_shading_rate_palettes              &ShadingRatePaletteNV
} 

// PhysicalDeviceShadingRateImageFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShadingRateImageFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shading_rate_image     Bool32
    shading_rate_coarse_sample_order Bool32
} 

// PhysicalDeviceShadingRateImagePropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceShadingRateImagePropertiesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shading_rate_texel_size Extent2D
    shading_rate_palette_size u32
    shading_rate_max_coarse_samples u32
} 

pub struct CoarseSampleLocationNV {
mut:
    pixel_x         u32
    pixel_y         u32
    sample          u32
} 

pub struct CoarseSampleOrderCustomNV {
mut:
    shading_rate                           ShadingRatePaletteEntryNV
    sample_count                           u32
    sample_location_count                  u32
    p_sample_locations                     &CoarseSampleLocationNV
} 

// PipelineViewportCoarseSampleOrderStateCreateInfoNV extends VkPipelineViewportStateCreateInfo
pub struct PipelineViewportCoarseSampleOrderStateCreateInfoNV {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    sample_order_type                         CoarseSampleOrderTypeNV
    custom_sample_order_count                 u32
    p_custom_sample_orders                    &CoarseSampleOrderCustomNV
} 

type VkCmdBindShadingRateImageNV = fn (     C.CommandBuffer,     C.ImageView,     ImageLayout) 

pub fn cmd_bind_shading_rate_image_nv(
    command_buffer                                  C.CommandBuffer,
    image_view                                      C.ImageView,
    image_layout                                    ImageLayout)  {
      f := VkCmdBindShadingRateImageNV((*loader_p).get_sym('vkCmdBindShadingRateImageNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindShadingRateImageNV': ${err}")
        return 
    })
    f(
    command_buffer,
    image_view,
    image_layout)
}


type VkCmdSetViewportShadingRatePaletteNV = fn (     C.CommandBuffer,     u32,     u32,     &ShadingRatePaletteNV) 

pub fn cmd_set_viewport_shading_rate_palette_nv(
    command_buffer                                  C.CommandBuffer,
    first_viewport                                  u32,
    viewport_count                                  u32,
    p_shading_rate_palettes                         &ShadingRatePaletteNV)  {
      f := VkCmdSetViewportShadingRatePaletteNV((*loader_p).get_sym('vkCmdSetViewportShadingRatePaletteNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetViewportShadingRatePaletteNV': ${err}")
        return 
    })
    f(
    command_buffer,
    first_viewport,
    viewport_count,
    p_shading_rate_palettes)
}


type VkCmdSetCoarseSampleOrderNV = fn (     C.CommandBuffer,     CoarseSampleOrderTypeNV,     u32,     &CoarseSampleOrderCustomNV) 

pub fn cmd_set_coarse_sample_order_nv(
    command_buffer                                  C.CommandBuffer,
    sample_order_type                               CoarseSampleOrderTypeNV,
    custom_sample_order_count                       u32,
    p_custom_sample_orders                          &CoarseSampleOrderCustomNV)  {
      f := VkCmdSetCoarseSampleOrderNV((*loader_p).get_sym('vkCmdSetCoarseSampleOrderNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetCoarseSampleOrderNV': ${err}")
        return 
    })
    f(
    command_buffer,
    sample_order_type,
    custom_sample_order_count,
    p_custom_sample_orders)
}




// VK_NV_ray_tracing is a preprocessor guard. Do not pass it to API calls.
const nv_ray_tracing = 1
pub type C.AccelerationStructureNV = voidptr
pub const nv_ray_tracing_spec_version       = 3
pub const nv_ray_tracing_extension_name     = "VK_NV_ray_tracing"
pub const shader_unused_khr                 = ~u32(0)
pub const shader_unused_nv                  = shader_unused_khr

pub enum RayTracingShaderGroupTypeKHR {
    ray_tracing_shader_group_type_general_khr = int(0)
    ray_tracing_shader_group_type_triangles_hit_group_khr = int(1)
    ray_tracing_shader_group_type_procedural_hit_group_khr = int(2)
    ray_tracing_shader_group_type_max_enum_khr = int(0x7FFFFFFF)
}

pub type RayTracingShaderGroupTypeNV = RayTracingShaderGroupTypeKHR


pub enum GeometryTypeKHR {
    geometry_type_triangles_khr = int(0)
    geometry_type_aabbs_khr = int(1)
    geometry_type_instances_khr = int(2)
    geometry_type_max_enum_khr = int(0x7FFFFFFF)
}

pub type GeometryTypeNV = GeometryTypeKHR


pub enum AccelerationStructureTypeKHR {
    acceleration_structure_type_top_level_khr = int(0)
    acceleration_structure_type_bottom_level_khr = int(1)
    acceleration_structure_type_generic_khr = int(2)
    acceleration_structure_type_max_enum_khr = int(0x7FFFFFFF)
}

pub type AccelerationStructureTypeNV = AccelerationStructureTypeKHR


pub enum CopyAccelerationStructureModeKHR {
    copy_acceleration_structure_mode_clone_khr = int(0)
    copy_acceleration_structure_mode_compact_khr = int(1)
    copy_acceleration_structure_mode_serialize_khr = int(2)
    copy_acceleration_structure_mode_deserialize_khr = int(3)
    copy_acceleration_structure_mode_max_enum_khr = int(0x7FFFFFFF)
}

pub type CopyAccelerationStructureModeNV = CopyAccelerationStructureModeKHR


pub enum AccelerationStructureMemoryRequirementsTypeNV {
    acceleration_structure_memory_requirements_type_object_nv = int(0)
    acceleration_structure_memory_requirements_type_build_scratch_nv = int(1)
    acceleration_structure_memory_requirements_type_update_scratch_nv = int(2)
    acceleration_structure_memory_requirements_type_max_enum_nv = int(0x7FFFFFFF)
}


pub enum GeometryFlagBitsKHR {
    geometry_opaque_bit_khr = int(0x00000001)
    geometry_no_duplicate_any_hit_invocation_bit_khr = int(0x00000002)
    geometry_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type GeometryFlagsKHR = u32
pub type GeometryFlagBitsNV = GeometryFlagBitsKHR


pub enum GeometryInstanceFlagBitsKHR {
    geometry_instance_triangle_facing_cull_disable_bit_khr = int(0x00000001)
    geometry_instance_triangle_flip_facing_bit_khr = int(0x00000002)
    geometry_instance_force_opaque_bit_khr = int(0x00000004)
    geometry_instance_force_no_opaque_bit_khr = int(0x00000008)
    geometry_instance_force_opacity_micromap_2_state_ext = int(0x00000010)
    geometry_instance_disable_opacity_micromaps_ext = int(0x00000020)
    geometry_instance_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type GeometryInstanceFlagsKHR = u32
pub type GeometryInstanceFlagBitsNV = GeometryInstanceFlagBitsKHR


pub enum BuildAccelerationStructureFlagBitsKHR {
    build_acceleration_structure_allow_update_bit_khr = int(0x00000001)
    build_acceleration_structure_allow_compaction_bit_khr = int(0x00000002)
    build_acceleration_structure_prefer_fast_trace_bit_khr = int(0x00000004)
    build_acceleration_structure_prefer_fast_build_bit_khr = int(0x00000008)
    build_acceleration_structure_low_memory_bit_khr = int(0x00000010)
    build_acceleration_structure_motion_bit_nv = int(0x00000020)
    build_acceleration_structure_allow_opacity_micromap_update_ext = int(0x00000040)
    build_acceleration_structure_allow_disable_opacity_micromaps_ext = int(0x00000080)
    build_acceleration_structure_allow_opacity_micromap_data_update_ext = int(0x00000100)
    build_acceleration_structure_allow_data_access_khr = int(0x00000800)
    build_acceleration_structure_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type BuildAccelerationStructureFlagsKHR = u32
pub type BuildAccelerationStructureFlagBitsNV = BuildAccelerationStructureFlagBitsKHR

pub struct RayTracingShaderGroupCreateInfoNV {
mut:
    s_type                                StructureType
    p_next                                voidptr
    vktype                                RayTracingShaderGroupTypeKHR
    general_shader                        u32
    closest_hit_shader                    u32
    any_hit_shader                        u32
    intersection_shader                   u32
} 

pub struct RayTracingPipelineCreateInfoNV {
mut:
    s_type                                            StructureType
    p_next                                            voidptr
    flags                                             PipelineCreateFlags
    stage_count                                       u32
    p_stages                                          &PipelineShaderStageCreateInfo
    group_count                                       u32
    p_groups                                          &RayTracingShaderGroupCreateInfoNV
    max_recursion_depth                               u32
    layout                                            C.PipelineLayout
    base_pipeline_handle                              C.Pipeline
    base_pipeline_index                               i32
} 

pub struct GeometryTrianglesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    vertex_data            C.Buffer
    vertex_offset          DeviceSize
    vertex_count           u32
    vertex_stride          DeviceSize
    vertex_format          Format
    index_data             C.Buffer
    index_offset           DeviceSize
    index_count            u32
    index_type             IndexType
    transform_data         C.Buffer
    transform_offset       DeviceSize
} 

pub struct GeometryAABBNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    aabb_data              C.Buffer
    num_aab_bs             u32
    stride                 u32
    offset                 DeviceSize
} 

pub struct GeometryDataNV {
mut:
    triangles                    GeometryTrianglesNV
    aabbs                        GeometryAABBNV
} 

pub struct GeometryNV {
mut:
    s_type                    StructureType
    p_next                    voidptr
    geometry_type             GeometryTypeKHR
    geometry                  GeometryDataNV
    flags                     GeometryFlagsKHR
} 

pub struct AccelerationStructureInfoNV {
mut:
    s_type                                     StructureType
    p_next                                     voidptr
    vktype                                     AccelerationStructureTypeNV
    flags                                      Flags
    instance_count                             u32
    geometry_count                             u32
    p_geometries                               &GeometryNV
} 

pub struct AccelerationStructureCreateInfoNV {
mut:
    s_type                               StructureType
    p_next                               voidptr
    compacted_size                       DeviceSize
    info                                 AccelerationStructureInfoNV
} 

pub struct BindAccelerationStructureMemoryInfoNV {
mut:
    s_type                           StructureType
    p_next                           voidptr
    acceleration_structure           C.AccelerationStructureNV
    memory                           C.DeviceMemory
    memory_offset                    DeviceSize
    device_index_count               u32
    p_device_indices                 &u32
} 

// WriteDescriptorSetAccelerationStructureNV extends VkWriteDescriptorSet
pub struct WriteDescriptorSetAccelerationStructureNV {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    acceleration_structure_count            u32
    p_acceleration_structures               &C.AccelerationStructureNV
} 

pub struct AccelerationStructureMemoryRequirementsInfoNV {
mut:
    s_type                                                 StructureType
    p_next                                                 voidptr
    vktype                                                 AccelerationStructureMemoryRequirementsTypeNV
    acceleration_structure                                 C.AccelerationStructureNV
} 

// PhysicalDeviceRayTracingPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceRayTracingPropertiesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_group_handle_size u32
    max_recursion_depth    u32
    max_shader_group_stride u32
    shader_group_base_alignment u32
    max_geometry_count     u64
    max_instance_count     u64
    max_triangle_count     u64
    max_descriptor_set_acceleration_structures u32
} 

pub struct TransformMatrixKHR {
mut:
    matrix[4]    []f32
} 

pub type TransformMatrixNV = TransformMatrixKHR

pub struct AabbPositionsKHR {
mut:
    min_x        f32
    min_y        f32
    min_z        f32
    max_x        f32
    max_y        f32
    max_z        f32
} 

pub type AabbPositionsNV = AabbPositionsKHR

pub struct AccelerationStructureInstanceKHR {
mut:
    transform                         TransformMatrixKHR
    instance_custom_index             u32
    mask                              u32
    instance_shader_binding_table_record_offset u32
    flags                             GeometryInstanceFlagsKHR
    acceleration_structure_reference  u64
} 

pub type AccelerationStructureInstanceNV = AccelerationStructureInstanceKHR

type VkCreateAccelerationStructureNV = fn (     C.Device,     &AccelerationStructureCreateInfoNV,     &AllocationCallbacks,     &C.AccelerationStructureNV) Result

pub fn create_acceleration_structure_nv(
    device                                          C.Device,
    p_create_info                                   &AccelerationStructureCreateInfoNV,
    p_allocator                                     &AllocationCallbacks,
    p_acceleration_structure                        &C.AccelerationStructureNV) Result {
      f := VkCreateAccelerationStructureNV((*loader_p).get_sym('vkCreateAccelerationStructureNV'
    ) or { 
        println("Couldn't load symbol for 'vkCreateAccelerationStructureNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_acceleration_structure)
}


type VkDestroyAccelerationStructureNV = fn (     C.Device,     C.AccelerationStructureNV,     &AllocationCallbacks) 

pub fn destroy_acceleration_structure_nv(
    device                                          C.Device,
    acceleration_structure                          C.AccelerationStructureNV,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyAccelerationStructureNV((*loader_p).get_sym('vkDestroyAccelerationStructureNV'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyAccelerationStructureNV': ${err}")
        return 
    })
    f(
    device,
    acceleration_structure,
    p_allocator)
}


type VkGetAccelerationStructureMemoryRequirementsNV = fn (     C.Device,     &AccelerationStructureMemoryRequirementsInfoNV,     &MemoryRequirements2KHR) 

pub fn get_acceleration_structure_memory_requirements_nv(
    device                                          C.Device,
    p_info                                          &AccelerationStructureMemoryRequirementsInfoNV,
    p_memory_requirements                           &MemoryRequirements2KHR)  {
      f := VkGetAccelerationStructureMemoryRequirementsNV((*loader_p).get_sym('vkGetAccelerationStructureMemoryRequirementsNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetAccelerationStructureMemoryRequirementsNV': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_memory_requirements)
}


type VkBindAccelerationStructureMemoryNV = fn (     C.Device,     u32,     &BindAccelerationStructureMemoryInfoNV) Result

pub fn bind_acceleration_structure_memory_nv(
    device                                          C.Device,
    bind_info_count                                 u32,
    p_bind_infos                                    &BindAccelerationStructureMemoryInfoNV) Result {
      f := VkBindAccelerationStructureMemoryNV((*loader_p).get_sym('vkBindAccelerationStructureMemoryNV'
    ) or { 
        println("Couldn't load symbol for 'vkBindAccelerationStructureMemoryNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    bind_info_count,
    p_bind_infos)
}


type VkCmdBuildAccelerationStructureNV = fn (     C.CommandBuffer,     &AccelerationStructureInfoNV,     C.Buffer,     DeviceSize,     Bool32,     C.AccelerationStructureNV,     C.AccelerationStructureNV,     C.Buffer,     DeviceSize) 

pub fn cmd_build_acceleration_structure_nv(
    command_buffer                                  C.CommandBuffer,
    p_info                                          &AccelerationStructureInfoNV,
    instance_data                                   C.Buffer,
    instance_offset                                 DeviceSize,
    update                                          Bool32,
    dst                                             C.AccelerationStructureNV,
    src                                             C.AccelerationStructureNV,
    scratch                                         C.Buffer,
    scratch_offset                                  DeviceSize)  {
      f := VkCmdBuildAccelerationStructureNV((*loader_p).get_sym('vkCmdBuildAccelerationStructureNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBuildAccelerationStructureNV': ${err}")
        return 
    })
    f(
    command_buffer,
    p_info,
    instance_data,
    instance_offset,
    update,
    dst,
    src,
    scratch,
    scratch_offset)
}


type VkCmdCopyAccelerationStructureNV = fn (     C.CommandBuffer,     C.AccelerationStructureNV,     C.AccelerationStructureNV,     CopyAccelerationStructureModeKHR) 

pub fn cmd_copy_acceleration_structure_nv(
    command_buffer                                  C.CommandBuffer,
    dst                                             C.AccelerationStructureNV,
    src                                             C.AccelerationStructureNV,
    mode                                            CopyAccelerationStructureModeKHR)  {
      f := VkCmdCopyAccelerationStructureNV((*loader_p).get_sym('vkCmdCopyAccelerationStructureNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyAccelerationStructureNV': ${err}")
        return 
    })
    f(
    command_buffer,
    dst,
    src,
    mode)
}


type VkCmdTraceRaysNV = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     C.Buffer,     DeviceSize,     DeviceSize,     C.Buffer,     DeviceSize,     DeviceSize,     C.Buffer,     DeviceSize,     DeviceSize,     u32,     u32,     u32) 

pub fn cmd_trace_rays_nv(
    command_buffer                                  C.CommandBuffer,
    raygen_shader_binding_table_buffer              C.Buffer,
    raygen_shader_binding_offset                    DeviceSize,
    miss_shader_binding_table_buffer                C.Buffer,
    miss_shader_binding_offset                      DeviceSize,
    miss_shader_binding_stride                      DeviceSize,
    hit_shader_binding_table_buffer                 C.Buffer,
    hit_shader_binding_offset                       DeviceSize,
    hit_shader_binding_stride                       DeviceSize,
    callable_shader_binding_table_buffer            C.Buffer,
    callable_shader_binding_offset                  DeviceSize,
    callable_shader_binding_stride                  DeviceSize,
    width                                           u32,
    height                                          u32,
    depth                                           u32)  {
      f := VkCmdTraceRaysNV((*loader_p).get_sym('vkCmdTraceRaysNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdTraceRaysNV': ${err}")
        return 
    })
    f(
    command_buffer,
    raygen_shader_binding_table_buffer,
    raygen_shader_binding_offset,
    miss_shader_binding_table_buffer,
    miss_shader_binding_offset,
    miss_shader_binding_stride,
    hit_shader_binding_table_buffer,
    hit_shader_binding_offset,
    hit_shader_binding_stride,
    callable_shader_binding_table_buffer,
    callable_shader_binding_offset,
    callable_shader_binding_stride,
    width,
    height,
    depth)
}


type VkCreateRayTracingPipelinesNV = fn (     C.Device,     C.PipelineCache,     u32,     &RayTracingPipelineCreateInfoNV,     &AllocationCallbacks,     &C.Pipeline) Result

pub fn create_ray_tracing_pipelines_nv(
    device                                          C.Device,
    pipeline_cache                                  C.PipelineCache,
    create_info_count                               u32,
    p_create_infos                                  &RayTracingPipelineCreateInfoNV,
    p_allocator                                     &AllocationCallbacks,
    p_pipelines                                     &C.Pipeline) Result {
      f := VkCreateRayTracingPipelinesNV((*loader_p).get_sym('vkCreateRayTracingPipelinesNV'
    ) or { 
        println("Couldn't load symbol for 'vkCreateRayTracingPipelinesNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    pipeline_cache,
    create_info_count,
    p_create_infos,
    p_allocator,
    p_pipelines)
}


type VkGetRayTracingShaderGroupHandlesKHR = fn (     C.Device,     C.Pipeline,     u32,     u32,     usize,     voidptr) Result

pub fn get_ray_tracing_shader_group_handles_khr(
    device                                          C.Device,
    pipeline                                        C.Pipeline,
    first_group                                     u32,
    group_count                                     u32,
    data_size                                       usize,
    p_data                                          voidptr) Result {
      f := VkGetRayTracingShaderGroupHandlesKHR((*loader_p).get_sym('vkGetRayTracingShaderGroupHandlesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetRayTracingShaderGroupHandlesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    pipeline,
    first_group,
    group_count,
    data_size,
    p_data)
}


type VkGetRayTracingShaderGroupHandlesNV = fn (     C.Device,     C.Pipeline,     u32,     u32,     usize,     voidptr) Result

pub fn get_ray_tracing_shader_group_handles_nv(
    device                                          C.Device,
    pipeline                                        C.Pipeline,
    first_group                                     u32,
    group_count                                     u32,
    data_size                                       usize,
    p_data                                          voidptr) Result {
      f := VkGetRayTracingShaderGroupHandlesNV((*loader_p).get_sym('vkGetRayTracingShaderGroupHandlesNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetRayTracingShaderGroupHandlesNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    pipeline,
    first_group,
    group_count,
    data_size,
    p_data)
}


type VkGetAccelerationStructureHandleNV = fn (     C.Device,     C.AccelerationStructureNV,     usize,     voidptr) Result

pub fn get_acceleration_structure_handle_nv(
    device                                          C.Device,
    acceleration_structure                          C.AccelerationStructureNV,
    data_size                                       usize,
    p_data                                          voidptr) Result {
      f := VkGetAccelerationStructureHandleNV((*loader_p).get_sym('vkGetAccelerationStructureHandleNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetAccelerationStructureHandleNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    acceleration_structure,
    data_size,
    p_data)
}


type VkCmdWriteAccelerationStructuresPropertiesNV = fn (     C.CommandBuffer,     u32,     &C.AccelerationStructureNV,     QueryType,     C.QueryPool,     u32) 

pub fn cmd_write_acceleration_structures_properties_nv(
    command_buffer                                  C.CommandBuffer,
    acceleration_structure_count                    u32,
    p_acceleration_structures                       &C.AccelerationStructureNV,
    query_type                                      QueryType,
    query_pool                                      C.QueryPool,
    first_query                                     u32)  {
      f := VkCmdWriteAccelerationStructuresPropertiesNV((*loader_p).get_sym('vkCmdWriteAccelerationStructuresPropertiesNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdWriteAccelerationStructuresPropertiesNV': ${err}")
        return 
    })
    f(
    command_buffer,
    acceleration_structure_count,
    p_acceleration_structures,
    query_type,
    query_pool,
    first_query)
}


type VkCompileDeferredNV = fn (     C.Device,     C.Pipeline,     u32) Result

pub fn compile_deferred_nv(
    device                                          C.Device,
    pipeline                                        C.Pipeline,
    shader                                          u32) Result {
      f := VkCompileDeferredNV((*loader_p).get_sym('vkCompileDeferredNV'
    ) or { 
        println("Couldn't load symbol for 'vkCompileDeferredNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    pipeline,
    shader)
}




// VK_NV_representative_fragment_test is a preprocessor guard. Do not pass it to API calls.
const nv_representative_fragment_test = 1
pub const nv_representative_fragment_test_spec_version = 2
pub const nv_representative_fragment_test_extension_name = "VK_NV_representative_fragment_test"
// PhysicalDeviceRepresentativeFragmentTestFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRepresentativeFragmentTestFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    representative_fragment_test Bool32
} 

// PipelineRepresentativeFragmentTestStateCreateInfoNV extends VkGraphicsPipelineCreateInfo
pub struct PipelineRepresentativeFragmentTestStateCreateInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    representative_fragment_test_enable Bool32
} 



// VK_EXT_filter_cubic is a preprocessor guard. Do not pass it to API calls.
const ext_filter_cubic = 1
pub const ext_filter_cubic_spec_version     = 3
pub const ext_filter_cubic_extension_name   = "VK_EXT_filter_cubic"
// PhysicalDeviceImageViewImageFormatInfoEXT extends VkPhysicalDeviceImageFormatInfo2
pub struct PhysicalDeviceImageViewImageFormatInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image_view_type        ImageViewType
} 

// FilterCubicImageViewImageFormatPropertiesEXT extends VkImageFormatProperties2
pub struct FilterCubicImageViewImageFormatPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    filter_cubic           Bool32
    filter_cubic_minmax    Bool32
} 



// VK_QCOM_render_pass_shader_resolve is a preprocessor guard. Do not pass it to API calls.
const qcom_render_pass_shader_resolve = 1
pub const qcom_render_pass_shader_resolve_spec_version = 4
pub const qcom_render_pass_shader_resolve_extension_name = "VK_QCOM_render_pass_shader_resolve"


// VK_EXT_global_priority is a preprocessor guard. Do not pass it to API calls.
const ext_global_priority = 1
pub const ext_global_priority_spec_version  = 2
pub const ext_global_priority_extension_name = "VK_EXT_global_priority"
pub type QueueGlobalPriorityEXT = QueueGlobalPriorityKHR

pub type DeviceQueueGlobalPriorityCreateInfoEXT = DeviceQueueGlobalPriorityCreateInfoKHR



// VK_EXT_external_memory_host is a preprocessor guard. Do not pass it to API calls.
const ext_external_memory_host = 1
pub const ext_external_memory_host_spec_version = 1
pub const ext_external_memory_host_extension_name = "VK_EXT_external_memory_host"
// ImportMemoryHostPointerInfoEXT extends VkMemoryAllocateInfo
pub struct ImportMemoryHostPointerInfoEXT {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    handle_type                               ExternalMemoryHandleTypeFlagBits
    p_host_pointer                            voidptr
} 

pub struct MemoryHostPointerPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    memory_type_bits       u32
} 

// PhysicalDeviceExternalMemoryHostPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceExternalMemoryHostPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    min_imported_host_pointer_alignment DeviceSize
} 

type VkGetMemoryHostPointerPropertiesEXT = fn (     C.Device,     ExternalMemoryHandleTypeFlagBits,     voidptr,     &MemoryHostPointerPropertiesEXT) Result

pub fn get_memory_host_pointer_properties_ext(
    device                                          C.Device,
    handle_type                                     ExternalMemoryHandleTypeFlagBits,
    p_host_pointer                                  voidptr,
    p_memory_host_pointer_properties                &MemoryHostPointerPropertiesEXT) Result {
      f := VkGetMemoryHostPointerPropertiesEXT((*loader_p).get_sym('vkGetMemoryHostPointerPropertiesEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetMemoryHostPointerPropertiesEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    handle_type,
    p_host_pointer,
    p_memory_host_pointer_properties)
}




// VK_AMD_buffer_marker is a preprocessor guard. Do not pass it to API calls.
const amd_buffer_marker = 1
pub const amd_buffer_marker_spec_version    = 1
pub const amd_buffer_marker_extension_name  = "VK_AMD_buffer_marker"
type VkCmdWriteBufferMarkerAMD = fn (     C.CommandBuffer,     PipelineStageFlagBits,     C.Buffer,     DeviceSize,     u32) 

pub fn cmd_write_buffer_marker_amd(
    command_buffer                                  C.CommandBuffer,
    pipeline_stage                                  PipelineStageFlagBits,
    dst_buffer                                      C.Buffer,
    dst_offset                                      DeviceSize,
    marker                                          u32)  {
      f := VkCmdWriteBufferMarkerAMD((*loader_p).get_sym('vkCmdWriteBufferMarkerAMD'
    ) or { 
        println("Couldn't load symbol for 'vkCmdWriteBufferMarkerAMD': ${err}")
        return 
    })
    f(
    command_buffer,
    pipeline_stage,
    dst_buffer,
    dst_offset,
    marker)
}




// VK_AMD_pipeline_compiler_control is a preprocessor guard. Do not pass it to API calls.
const amd_pipeline_compiler_control = 1
pub const amd_pipeline_compiler_control_spec_version = 1
pub const amd_pipeline_compiler_control_extension_name = "VK_AMD_pipeline_compiler_control"

pub enum PipelineCompilerControlFlagBitsAMD {
    pipeline_compiler_control_flag_bits_max_enum_amd = int(0x7FFFFFFF)
}

pub type PipelineCompilerControlFlagsAMD = u32
// PipelineCompilerControlCreateInfoAMD extends VkGraphicsPipelineCreateInfo,VkComputePipelineCreateInfo,VkExecutionGraphPipelineCreateInfoAMDX
pub struct PipelineCompilerControlCreateInfoAMD {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    compiler_control_flags                   PipelineCompilerControlFlagsAMD
} 



// VK_EXT_calibrated_timestamps is a preprocessor guard. Do not pass it to API calls.
const ext_calibrated_timestamps = 1
pub const ext_calibrated_timestamps_spec_version = 2
pub const ext_calibrated_timestamps_extension_name = "VK_EXT_calibrated_timestamps"

pub enum TimeDomainEXT {
    time_domain_device_ext = int(0)
    time_domain_clock_monotonic_ext = int(1)
    time_domain_clock_monotonic_raw_ext = int(2)
    time_domain_query_performance_counter_ext = int(3)
    time_domain_max_enum_ext = int(0x7FFFFFFF)
}

pub struct CalibratedTimestampInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    time_domain            TimeDomainEXT
} 

type VkGetPhysicalDeviceCalibrateableTimeDomainsEXT = fn (     C.PhysicalDevice,     &u32,     &TimeDomainEXT) Result

pub fn get_physical_device_calibrateable_time_domains_ext(
    physical_device                                 C.PhysicalDevice,
    p_time_domain_count                             &u32,
    p_time_domains                                  &TimeDomainEXT) Result {
      f := VkGetPhysicalDeviceCalibrateableTimeDomainsEXT((*loader_p).get_sym('vkGetPhysicalDeviceCalibrateableTimeDomainsEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceCalibrateableTimeDomainsEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_time_domain_count,
    p_time_domains)
}


type VkGetCalibratedTimestampsEXT = fn (     C.Device,     u32,     &CalibratedTimestampInfoEXT,     &u64,     &u64) Result

pub fn get_calibrated_timestamps_ext(
    device                                          C.Device,
    timestamp_count                                 u32,
    p_timestamp_infos                               &CalibratedTimestampInfoEXT,
    p_timestamps                                    &u64,
    p_max_deviation                                 &u64) Result {
      f := VkGetCalibratedTimestampsEXT((*loader_p).get_sym('vkGetCalibratedTimestampsEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetCalibratedTimestampsEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    timestamp_count,
    p_timestamp_infos,
    p_timestamps,
    p_max_deviation)
}




// VK_AMD_shader_core_properties is a preprocessor guard. Do not pass it to API calls.
const amd_shader_core_properties = 1
pub const amd_shader_core_properties_spec_version = 2
pub const amd_shader_core_properties_extension_name = "VK_AMD_shader_core_properties"
// PhysicalDeviceShaderCorePropertiesAMD extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceShaderCorePropertiesAMD {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_engine_count    u32
    shader_arrays_per_engine_count u32
    compute_units_per_shader_array u32
    simd_per_compute_unit  u32
    wavefronts_per_simd    u32
    wavefront_size         u32
    sgprs_per_simd         u32
    min_sgpr_allocation    u32
    max_sgpr_allocation    u32
    sgpr_allocation_granularity u32
    vgprs_per_simd         u32
    min_vgpr_allocation    u32
    max_vgpr_allocation    u32
    vgpr_allocation_granularity u32
} 



// VK_AMD_memory_overallocation_behavior is a preprocessor guard. Do not pass it to API calls.
const amd_memory_overallocation_behavior = 1
pub const amd_memory_overallocation_behavior_spec_version = 1
pub const amd_memory_overallocation_behavior_extension_name = "VK_AMD_memory_overallocation_behavior"

pub enum MemoryOverallocationBehaviorAMD {
    memory_overallocation_behavior_default_amd = int(0)
    memory_overallocation_behavior_allowed_amd = int(1)
    memory_overallocation_behavior_disallowed_amd = int(2)
    memory_overallocation_behavior_max_enum_amd = int(0x7FFFFFFF)
}

// DeviceMemoryOverallocationCreateInfoAMD extends VkDeviceCreateInfo
pub struct DeviceMemoryOverallocationCreateInfoAMD {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    overallocation_behavior                  MemoryOverallocationBehaviorAMD
} 



// VK_EXT_vertex_attribute_divisor is a preprocessor guard. Do not pass it to API calls.
const ext_vertex_attribute_divisor = 1
pub const ext_vertex_attribute_divisor_spec_version = 3
pub const ext_vertex_attribute_divisor_extension_name = "VK_EXT_vertex_attribute_divisor"
// PhysicalDeviceVertexAttributeDivisorPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceVertexAttributeDivisorPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_vertex_attrib_divisor u32
} 

pub struct VertexInputBindingDivisorDescriptionEXT {
mut:
    binding         u32
    divisor         u32
} 

// PipelineVertexInputDivisorStateCreateInfoEXT extends VkPipelineVertexInputStateCreateInfo
pub struct PipelineVertexInputDivisorStateCreateInfoEXT {
mut:
    s_type                                                  StructureType
    p_next                                                  voidptr
    vertex_binding_divisor_count                            u32
    p_vertex_binding_divisors                               &VertexInputBindingDivisorDescriptionEXT
} 

// PhysicalDeviceVertexAttributeDivisorFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceVertexAttributeDivisorFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    vertex_attribute_instance_rate_divisor Bool32
    vertex_attribute_instance_rate_zero_divisor Bool32
} 



// VK_GGP_frame_token is a preprocessor guard. Do not pass it to API calls.
const ggp_frame_token = 1
pub const ggp_frame_token_spec_version      = 1
pub const ggp_frame_token_extension_name    = "VK_GGP_frame_token"
// PresentFrameTokenGGP extends VkPresentInfoKHR
pub struct PresentFrameTokenGGP {
mut:
    s_type                 StructureType
    p_next                 voidptr
    frame_token            u64
} 



// VK_EXT_pipeline_creation_feedback is a preprocessor guard. Do not pass it to API calls.
const ext_pipeline_creation_feedback = 1
pub const ext_pipeline_creation_feedback_spec_version = 1
pub const ext_pipeline_creation_feedback_extension_name = "VK_EXT_pipeline_creation_feedback"
pub type PipelineCreationFeedbackFlagBitsEXT = PipelineCreationFeedbackFlagBits

pub type PipelineCreationFeedbackCreateInfoEXT = PipelineCreationFeedbackCreateInfo

pub type PipelineCreationFeedbackEXT = PipelineCreationFeedback



// VK_NV_shader_subgroup_partitioned is a preprocessor guard. Do not pass it to API calls.
const nv_shader_subgroup_partitioned = 1
pub const nv_shader_subgroup_partitioned_spec_version = 1
pub const nv_shader_subgroup_partitioned_extension_name = "VK_NV_shader_subgroup_partitioned"


// VK_NV_compute_shader_derivatives is a preprocessor guard. Do not pass it to API calls.
const nv_compute_shader_derivatives = 1
pub const nv_compute_shader_derivatives_spec_version = 1
pub const nv_compute_shader_derivatives_extension_name = "VK_NV_compute_shader_derivatives"
// PhysicalDeviceComputeShaderDerivativesFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceComputeShaderDerivativesFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    compute_derivative_group_quads Bool32
    compute_derivative_group_linear Bool32
} 



// VK_NV_mesh_shader is a preprocessor guard. Do not pass it to API calls.
const nv_mesh_shader = 1
pub const nv_mesh_shader_spec_version       = 1
pub const nv_mesh_shader_extension_name     = "VK_NV_mesh_shader"
// PhysicalDeviceMeshShaderFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMeshShaderFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    task_shader            Bool32
    mesh_shader            Bool32
} 

// PhysicalDeviceMeshShaderPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceMeshShaderPropertiesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_draw_mesh_tasks_count u32
    max_task_work_group_invocations u32
    max_task_work_group_size []u32
    max_task_total_memory_size u32
    max_task_output_count  u32
    max_mesh_work_group_invocations u32
    max_mesh_work_group_size []u32
    max_mesh_total_memory_size u32
    max_mesh_output_vertices u32
    max_mesh_output_primitives u32
    max_mesh_multiview_view_count u32
    mesh_output_per_vertex_granularity u32
    mesh_output_per_primitive_granularity u32
} 

pub struct DrawMeshTasksIndirectCommandNV {
mut:
    task_count      u32
    first_task      u32
} 

type VkCmdDrawMeshTasksNV = fn (     C.CommandBuffer,     u32,     u32) 

pub fn cmd_draw_mesh_tasks_nv(
    command_buffer                                  C.CommandBuffer,
    task_count                                      u32,
    first_task                                      u32)  {
      f := VkCmdDrawMeshTasksNV((*loader_p).get_sym('vkCmdDrawMeshTasksNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawMeshTasksNV': ${err}")
        return 
    })
    f(
    command_buffer,
    task_count,
    first_task)
}


type VkCmdDrawMeshTasksIndirectNV = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_mesh_tasks_indirect_nv(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    draw_count                                      u32,
    stride                                          u32)  {
      f := VkCmdDrawMeshTasksIndirectNV((*loader_p).get_sym('vkCmdDrawMeshTasksIndirectNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawMeshTasksIndirectNV': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    draw_count,
    stride)
}


type VkCmdDrawMeshTasksIndirectCountNV = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_mesh_tasks_indirect_count_nv(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    count_buffer                                    C.Buffer,
    count_buffer_offset                             DeviceSize,
    max_draw_count                                  u32,
    stride                                          u32)  {
      f := VkCmdDrawMeshTasksIndirectCountNV((*loader_p).get_sym('vkCmdDrawMeshTasksIndirectCountNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawMeshTasksIndirectCountNV': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    count_buffer,
    count_buffer_offset,
    max_draw_count,
    stride)
}




// VK_NV_fragment_shader_barycentric is a preprocessor guard. Do not pass it to API calls.
const nv_fragment_shader_barycentric = 1
pub const nv_fragment_shader_barycentric_spec_version = 1
pub const nv_fragment_shader_barycentric_extension_name = "VK_NV_fragment_shader_barycentric"
pub type PhysicalDeviceFragmentShaderBarycentricFeaturesNV = PhysicalDeviceFragmentShaderBarycentricFeaturesKHR



// VK_NV_shader_image_footprint is a preprocessor guard. Do not pass it to API calls.
const nv_shader_image_footprint = 1
pub const nv_shader_image_footprint_spec_version = 2
pub const nv_shader_image_footprint_extension_name = "VK_NV_shader_image_footprint"
// PhysicalDeviceShaderImageFootprintFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderImageFootprintFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image_footprint        Bool32
} 



// VK_NV_scissor_exclusive is a preprocessor guard. Do not pass it to API calls.
const nv_scissor_exclusive = 1
pub const nv_scissor_exclusive_spec_version = 2
pub const nv_scissor_exclusive_extension_name = "VK_NV_scissor_exclusive"
// PipelineViewportExclusiveScissorStateCreateInfoNV extends VkPipelineViewportStateCreateInfo
pub struct PipelineViewportExclusiveScissorStateCreateInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    exclusive_scissor_count u32
    p_exclusive_scissors   &Rect2D
} 

// PhysicalDeviceExclusiveScissorFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceExclusiveScissorFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    exclusive_scissor      Bool32
} 

type VkCmdSetExclusiveScissorEnableNV = fn (     C.CommandBuffer,     u32,     u32,     &Bool32) 

pub fn cmd_set_exclusive_scissor_enable_nv(
    command_buffer                                  C.CommandBuffer,
    first_exclusive_scissor                         u32,
    exclusive_scissor_count                         u32,
    p_exclusive_scissor_enables                     &Bool32)  {
      f := VkCmdSetExclusiveScissorEnableNV((*loader_p).get_sym('vkCmdSetExclusiveScissorEnableNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetExclusiveScissorEnableNV': ${err}")
        return 
    })
    f(
    command_buffer,
    first_exclusive_scissor,
    exclusive_scissor_count,
    p_exclusive_scissor_enables)
}


type VkCmdSetExclusiveScissorNV = fn (     C.CommandBuffer,     u32,     u32,     &Rect2D) 

pub fn cmd_set_exclusive_scissor_nv(
    command_buffer                                  C.CommandBuffer,
    first_exclusive_scissor                         u32,
    exclusive_scissor_count                         u32,
    p_exclusive_scissors                            &Rect2D)  {
      f := VkCmdSetExclusiveScissorNV((*loader_p).get_sym('vkCmdSetExclusiveScissorNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetExclusiveScissorNV': ${err}")
        return 
    })
    f(
    command_buffer,
    first_exclusive_scissor,
    exclusive_scissor_count,
    p_exclusive_scissors)
}




// VK_NV_device_diagnostic_checkpoints is a preprocessor guard. Do not pass it to API calls.
const nv_device_diagnostic_checkpoints = 1
pub const nv_device_diagnostic_checkpoints_spec_version = 2
pub const nv_device_diagnostic_checkpoints_extension_name = "VK_NV_device_diagnostic_checkpoints"
// QueueFamilyCheckpointPropertiesNV extends VkQueueFamilyProperties2
pub struct QueueFamilyCheckpointPropertiesNV {
mut:
    s_type                      StructureType
    p_next                      voidptr
    checkpoint_execution_stage_mask PipelineStageFlags
} 

pub struct CheckpointDataNV {
mut:
    s_type                         StructureType
    p_next                         voidptr
    stage                          PipelineStageFlagBits
    p_checkpoint_marker            voidptr
} 

type VkCmdSetCheckpointNV = fn (     C.CommandBuffer,     voidptr) 

pub fn cmd_set_checkpoint_nv(
    command_buffer                                  C.CommandBuffer,
    p_checkpoint_marker                             voidptr)  {
      f := VkCmdSetCheckpointNV((*loader_p).get_sym('vkCmdSetCheckpointNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetCheckpointNV': ${err}")
        return 
    })
    f(
    command_buffer,
    p_checkpoint_marker)
}


type VkGetQueueCheckpointDataNV = fn (     C.Queue,     &u32,     &CheckpointDataNV) 

pub fn get_queue_checkpoint_data_nv(
    queue                                           C.Queue,
    p_checkpoint_data_count                         &u32,
    p_checkpoint_data                               &CheckpointDataNV)  {
      f := VkGetQueueCheckpointDataNV((*loader_p).get_sym('vkGetQueueCheckpointDataNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetQueueCheckpointDataNV': ${err}")
        return 
    })
    f(
    queue,
    p_checkpoint_data_count,
    p_checkpoint_data)
}




// VK_INTEL_shader_integer_functions2 is a preprocessor guard. Do not pass it to API calls.
const intel_shader_integer_functions2 = 1
pub const intel_shader_integer_functions_2_spec_version = 1
pub const intel_shader_integer_functions_2_extension_name = "VK_INTE_shader_integer_functions2"
// PhysicalDeviceShaderIntegerFunctions2FeaturesINTEL extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderIntegerFunctions2FeaturesINTEL {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_integer_functions2 Bool32
} 



// VK_INTEL_performance_query is a preprocessor guard. Do not pass it to API calls.
const intel_performance_query = 1
pub type C.PerformanceConfigurationINTEL = voidptr
pub const intel_performance_query_spec_version = 2
pub const intel_performance_query_extension_name = "VK_INTE_performance_query"

pub enum PerformanceConfigurationTypeINTEL {
    performance_configuration_type_command_queue_metrics_discovery_activated_intel = int(0)
    performance_configuration_type_max_enum_intel = int(0x7FFFFFFF)
}


pub enum QueryPoolSamplingModeINTEL {
    query_pool_sampling_mode_manual_intel = int(0)
    query_pool_sampling_mode_max_enum_intel = int(0x7FFFFFFF)
}


pub enum PerformanceOverrideTypeINTEL {
    performance_override_type_null_hardware_intel = int(0)
    performance_override_type_flush_gpu_caches_intel = int(1)
    performance_override_type_max_enum_intel = int(0x7FFFFFFF)
}


pub enum PerformanceParameterTypeINTEL {
    performance_parameter_type_hw_counters_supported_intel = int(0)
    performance_parameter_type_stream_marker_valid_bits_intel = int(1)
    performance_parameter_type_max_enum_intel = int(0x7FFFFFFF)
}


pub enum PerformanceValueTypeINTEL {
    performance_value_type_uint32_intel = int(0)
    performance_value_type_uint64_intel = int(1)
    performance_value_type_float_intel = int(2)
    performance_value_type_bool_intel = int(3)
    performance_value_type_string_intel = int(4)
    performance_value_type_max_enum_intel = int(0x7FFFFFFF)
}

pub union PerformanceValueDataINTEL {
mut:
    value32            u32
    value64            u64
    value_float        f32
    value_bool         Bool32
    value_string       &char
} 

pub struct PerformanceValueINTEL {
mut:
    vktype                             PerformanceValueTypeINTEL
    data                               PerformanceValueDataINTEL
} 

pub struct InitializePerformanceApiInfoINTEL {
mut:
    s_type                 StructureType
    p_next                 voidptr
    p_user_data            voidptr
} 

// QueryPoolPerformanceQueryCreateInfoINTEL extends VkQueryPoolCreateInfo
pub struct QueryPoolPerformanceQueryCreateInfoINTEL {
mut:
    s_type                              StructureType
    p_next                              voidptr
    performance_counters_sampling       QueryPoolSamplingModeINTEL
} 

pub type QueryPoolCreateInfoINTEL = QueryPoolPerformanceQueryCreateInfoINTEL

pub struct PerformanceMarkerInfoINTEL {
mut:
    s_type                 StructureType
    p_next                 voidptr
    marker                 u64
} 

pub struct PerformanceStreamMarkerInfoINTEL {
mut:
    s_type                 StructureType
    p_next                 voidptr
    marker                 u32
} 

pub struct PerformanceOverrideInfoINTEL {
mut:
    s_type                                StructureType
    p_next                                voidptr
    vktype                                PerformanceOverrideTypeINTEL
    enable                                Bool32
    parameter                             u64
} 

pub struct PerformanceConfigurationAcquireInfoINTEL {
mut:
    s_type                                     StructureType
    p_next                                     voidptr
    vktype                                     PerformanceConfigurationTypeINTEL
} 

type VkInitializePerformanceApiINTEL = fn (     C.Device,     &InitializePerformanceApiInfoINTEL) Result

pub fn initialize_performance_api_intel(
    device                                          C.Device,
    p_initialize_info                               &InitializePerformanceApiInfoINTEL) Result {
      f := VkInitializePerformanceApiINTEL((*loader_p).get_sym('vkInitializePerformanceApiINTEL'
    ) or { 
        println("Couldn't load symbol for 'vkInitializePerformanceApiINTEL': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_initialize_info)
}


type VkUninitializePerformanceApiINTEL = fn (     C.Device) 

pub fn uninitialize_performance_api_intel(
    device                                          C.Device)  {
      f := VkUninitializePerformanceApiINTEL((*loader_p).get_sym('vkUninitializePerformanceApiINTEL'
    ) or { 
        println("Couldn't load symbol for 'vkUninitializePerformanceApiINTEL': ${err}")
        return 
    })
    f(
    device)
}


type VkCmdSetPerformanceMarkerINTEL = fn (     C.CommandBuffer,     &PerformanceMarkerInfoINTEL) Result

pub fn cmd_set_performance_marker_intel(
    command_buffer                                  C.CommandBuffer,
    p_marker_info                                   &PerformanceMarkerInfoINTEL) Result {
      f := VkCmdSetPerformanceMarkerINTEL((*loader_p).get_sym('vkCmdSetPerformanceMarkerINTEL'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetPerformanceMarkerINTEL': ${err}")
        return Result.error_unknown
    })
    return f(
    command_buffer,
    p_marker_info)
}


type VkCmdSetPerformanceStreamMarkerINTEL = fn (     C.CommandBuffer,     &PerformanceStreamMarkerInfoINTEL) Result

pub fn cmd_set_performance_stream_marker_intel(
    command_buffer                                  C.CommandBuffer,
    p_marker_info                                   &PerformanceStreamMarkerInfoINTEL) Result {
      f := VkCmdSetPerformanceStreamMarkerINTEL((*loader_p).get_sym('vkCmdSetPerformanceStreamMarkerINTEL'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetPerformanceStreamMarkerINTEL': ${err}")
        return Result.error_unknown
    })
    return f(
    command_buffer,
    p_marker_info)
}


type VkCmdSetPerformanceOverrideINTEL = fn (     C.CommandBuffer,     &PerformanceOverrideInfoINTEL) Result

pub fn cmd_set_performance_override_intel(
    command_buffer                                  C.CommandBuffer,
    p_override_info                                 &PerformanceOverrideInfoINTEL) Result {
      f := VkCmdSetPerformanceOverrideINTEL((*loader_p).get_sym('vkCmdSetPerformanceOverrideINTEL'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetPerformanceOverrideINTEL': ${err}")
        return Result.error_unknown
    })
    return f(
    command_buffer,
    p_override_info)
}


type VkAcquirePerformanceConfigurationINTEL = fn (     C.Device,     &PerformanceConfigurationAcquireInfoINTEL,     &C.PerformanceConfigurationINTEL) Result

pub fn acquire_performance_configuration_intel(
    device                                          C.Device,
    p_acquire_info                                  &PerformanceConfigurationAcquireInfoINTEL,
    p_configuration                                 &C.PerformanceConfigurationINTEL) Result {
      f := VkAcquirePerformanceConfigurationINTEL((*loader_p).get_sym('vkAcquirePerformanceConfigurationINTEL'
    ) or { 
        println("Couldn't load symbol for 'vkAcquirePerformanceConfigurationINTEL': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_acquire_info,
    p_configuration)
}


type VkReleasePerformanceConfigurationINTEL = fn (     C.Device,     C.PerformanceConfigurationINTEL) Result

pub fn release_performance_configuration_intel(
    device                                          C.Device,
    configuration                                   C.PerformanceConfigurationINTEL) Result {
      f := VkReleasePerformanceConfigurationINTEL((*loader_p).get_sym('vkReleasePerformanceConfigurationINTEL'
    ) or { 
        println("Couldn't load symbol for 'vkReleasePerformanceConfigurationINTEL': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    configuration)
}


type VkQueueSetPerformanceConfigurationINTEL = fn (     C.Queue,     C.PerformanceConfigurationINTEL) Result

pub fn queue_set_performance_configuration_intel(
    queue                                           C.Queue,
    configuration                                   C.PerformanceConfigurationINTEL) Result {
      f := VkQueueSetPerformanceConfigurationINTEL((*loader_p).get_sym('vkQueueSetPerformanceConfigurationINTEL'
    ) or { 
        println("Couldn't load symbol for 'vkQueueSetPerformanceConfigurationINTEL': ${err}")
        return Result.error_unknown
    })
    return f(
    queue,
    configuration)
}


type VkGetPerformanceParameterINTEL = fn (     C.Device,     PerformanceParameterTypeINTEL,     &PerformanceValueINTEL) Result

pub fn get_performance_parameter_intel(
    device                                          C.Device,
    parameter                                       PerformanceParameterTypeINTEL,
    p_value                                         &PerformanceValueINTEL) Result {
      f := VkGetPerformanceParameterINTEL((*loader_p).get_sym('vkGetPerformanceParameterINTEL'
    ) or { 
        println("Couldn't load symbol for 'vkGetPerformanceParameterINTEL': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    parameter,
    p_value)
}




// VK_EXT_pci_bus_info is a preprocessor guard. Do not pass it to API calls.
const ext_pci_bus_info = 1
pub const ext_pci_bus_info_spec_version     = 2
pub const ext_pci_bus_info_extension_name   = "VK_EXT_pci_bus_info"
// PhysicalDevicePCIBusInfoPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDevicePCIBusInfoPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pci_domain             u32
    pci_bus                u32
    pci_device             u32
    pci_function           u32
} 



// VK_AMD_display_native_hdr is a preprocessor guard. Do not pass it to API calls.
const amd_display_native_hdr = 1
pub const amd_display_native_hdr_spec_version = 1
pub const amd_display_native_hdr_extension_name = "VK_AMD_display_native_hdr"
// DisplayNativeHdrSurfaceCapabilitiesAMD extends VkSurfaceCapabilities2KHR
pub struct DisplayNativeHdrSurfaceCapabilitiesAMD {
mut:
    s_type                 StructureType
    p_next                 voidptr
    local_dimming_support  Bool32
} 

// SwapchainDisplayNativeHdrCreateInfoAMD extends VkSwapchainCreateInfoKHR
pub struct SwapchainDisplayNativeHdrCreateInfoAMD {
mut:
    s_type                 StructureType
    p_next                 voidptr
    local_dimming_enable   Bool32
} 

type VkSetLocalDimmingAMD = fn (     C.Device,     C.SwapchainKHR,     Bool32) 

pub fn set_local_dimming_amd(
    device                                          C.Device,
    swap_chain                                      C.SwapchainKHR,
    local_dimming_enable                            Bool32)  {
      f := VkSetLocalDimmingAMD((*loader_p).get_sym('vkSetLocalDimmingAMD'
    ) or { 
        println("Couldn't load symbol for 'vkSetLocalDimmingAMD': ${err}")
        return 
    })
    f(
    device,
    swap_chain,
    local_dimming_enable)
}




// VK_FUCHSIA_imagepipe_surface is a preprocessor guard. Do not pass it to API calls.
const fuchsia_imagepipe_surface = 1
pub const fuchsia_imagepipe_surface_spec_version = 1
pub const fuchsia_imagepipe_surface_extension_name = "VK_CHSIA_imagepipe_surface"
pub type ImagePipeSurfaceCreateFlagsFUCHSIA = u32
pub struct ImagePipeSurfaceCreateInfoFUCHSIA {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    flags                                       ImagePipeSurfaceCreateFlagsFUCHSIA
    image_pipe_handle                           voidptr
} 

type VkCreateImagePipeSurfaceFUCHSIA = fn (     C.Instance,     &ImagePipeSurfaceCreateInfoFUCHSIA,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_image_pipe_surface_fuchsia(
    instance                                        C.Instance,
    p_create_info                                   &ImagePipeSurfaceCreateInfoFUCHSIA,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateImagePipeSurfaceFUCHSIA((*loader_p).get_sym('vkCreateImagePipeSurfaceFUCHSIA'
    ) or { 
        println("Couldn't load symbol for 'vkCreateImagePipeSurfaceFUCHSIA': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}




// VK_EXT_metal_surface is a preprocessor guard. Do not pass it to API calls.
const ext_metal_surface = 1
pub const ext_metal_surface_spec_version    = 1
pub const ext_metal_surface_extension_name  = "VK_EXT_metal_surface"
pub type MetalSurfaceCreateFlagsEXT = u32
pub struct MetalSurfaceCreateInfoEXT {
mut:
    s_type                              StructureType
    p_next                              voidptr
    flags                               MetalSurfaceCreateFlagsEXT
    p_layer                             voidptr
} 

type VkCreateMetalSurfaceEXT = fn (     C.Instance,     &MetalSurfaceCreateInfoEXT,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_metal_surface_ext(
    instance                                        C.Instance,
    p_create_info                                   &MetalSurfaceCreateInfoEXT,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateMetalSurfaceEXT((*loader_p).get_sym('vkCreateMetalSurfaceEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCreateMetalSurfaceEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}




// VK_EXT_fragment_density_map is a preprocessor guard. Do not pass it to API calls.
const ext_fragment_density_map = 1
pub const ext_fragment_density_map_spec_version = 2
pub const ext_fragment_density_map_extension_name = "VK_EXT_fragment_density_map"
// PhysicalDeviceFragmentDensityMapFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceFragmentDensityMapFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    fragment_density_map   Bool32
    fragment_density_map_dynamic Bool32
    fragment_density_map_non_subsampled_images Bool32
} 

// PhysicalDeviceFragmentDensityMapPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceFragmentDensityMapPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    min_fragment_density_texel_size Extent2D
    max_fragment_density_texel_size Extent2D
    fragment_density_invocations Bool32
} 

// RenderPassFragmentDensityMapCreateInfoEXT extends VkRenderPassCreateInfo,VkRenderPassCreateInfo2
pub struct RenderPassFragmentDensityMapCreateInfoEXT {
mut:
    s_type                       StructureType
    p_next                       voidptr
    fragment_density_map_attachment AttachmentReference
} 



// VK_EXT_scalar_block_layout is a preprocessor guard. Do not pass it to API calls.
const ext_scalar_block_layout = 1
pub const ext_scalar_block_layout_spec_version = 1
pub const ext_scalar_block_layout_extension_name = "VK_EXT_scalar_block_layout"
pub type PhysicalDeviceScalarBlockLayoutFeaturesEXT = PhysicalDeviceScalarBlockLayoutFeatures



// VK_GOOGLE_hlsl_functionality1 is a preprocessor guard. Do not pass it to API calls.
const google_hlsl_functionality1 = 1
pub const google_hlsl_functionality_1_spec_version = 1
pub const google_hlsl_functionality_1_extension_name = "VK_GOOGE_hlsl_functionality1"
pub const google_hlsl_functionality1_spec_version = google_hlsl_functionality_1_spec_version
pub const google_hlsl_functionality1_extension_name = google_hlsl_functionality_1_extension_name


// VK_GOOGLE_decorate_string is a preprocessor guard. Do not pass it to API calls.
const google_decorate_string = 1
pub const google_decorate_string_spec_version = 1
pub const google_decorate_string_extension_name = "VK_GOOGE_decorate_string"


// VK_EXT_subgroup_size_control is a preprocessor guard. Do not pass it to API calls.
const ext_subgroup_size_control = 1
pub const ext_subgroup_size_control_spec_version = 2
pub const ext_subgroup_size_control_extension_name = "VK_EXT_subgroup_size_control"
pub type PhysicalDeviceSubgroupSizeControlFeaturesEXT = PhysicalDeviceSubgroupSizeControlFeatures

pub type PhysicalDeviceSubgroupSizeControlPropertiesEXT = PhysicalDeviceSubgroupSizeControlProperties

pub type PipelineShaderStageRequiredSubgroupSizeCreateInfoEXT = PipelineShaderStageRequiredSubgroupSizeCreateInfo



// VK_AMD_shader_core_properties2 is a preprocessor guard. Do not pass it to API calls.
const amd_shader_core_properties2 = 1
pub const amd_shader_core_properties_2_spec_version = 1
pub const amd_shader_core_properties_2_extension_name = "VK_AMD_shader_core_properties2"

pub enum ShaderCorePropertiesFlagBitsAMD {
    shader_core_properties_flag_bits_max_enum_amd = int(0x7FFFFFFF)
}

pub type ShaderCorePropertiesFlagsAMD = u32
// PhysicalDeviceShaderCoreProperties2AMD extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceShaderCoreProperties2AMD {
mut:
    s_type                                StructureType
    p_next                                voidptr
    shader_core_features                  ShaderCorePropertiesFlagsAMD
    active_compute_unit_count             u32
} 



// VK_AMD_device_coherent_memory is a preprocessor guard. Do not pass it to API calls.
const amd_device_coherent_memory = 1
pub const amd_device_coherent_memory_spec_version = 1
pub const amd_device_coherent_memory_extension_name = "VK_AMD_device_coherent_memory"
// PhysicalDeviceCoherentMemoryFeaturesAMD extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceCoherentMemoryFeaturesAMD {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_coherent_memory Bool32
} 



// VK_EXT_shader_image_atomic_int64 is a preprocessor guard. Do not pass it to API calls.
const ext_shader_image_atomic_int64 = 1
pub const ext_shader_image_atomic_int64_spec_version = 1
pub const ext_shader_image_atomic_int64_extension_name = "VK_EXT_shader_image_atomic_int64"
// PhysicalDeviceShaderImageAtomicInt64FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderImageAtomicInt64FeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_image_int64_atomics Bool32
    sparse_image_int64_atomics Bool32
} 



// VK_EXT_memory_budget is a preprocessor guard. Do not pass it to API calls.
const ext_memory_budget = 1
pub const ext_memory_budget_spec_version    = 1
pub const ext_memory_budget_extension_name  = "VK_EXT_memory_budget"
// PhysicalDeviceMemoryBudgetPropertiesEXT extends VkPhysicalDeviceMemoryProperties2
pub struct PhysicalDeviceMemoryBudgetPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    heap_budget            []DeviceSize
    heap_usage             []DeviceSize
} 



// VK_EXT_memory_priority is a preprocessor guard. Do not pass it to API calls.
const ext_memory_priority = 1
pub const ext_memory_priority_spec_version  = 1
pub const ext_memory_priority_extension_name = "VK_EXT_memory_priority"
// PhysicalDeviceMemoryPriorityFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMemoryPriorityFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    memory_priority        Bool32
} 

// MemoryPriorityAllocateInfoEXT extends VkMemoryAllocateInfo
pub struct MemoryPriorityAllocateInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    priority               f32
} 



// VK_NV_dedicated_allocation_image_aliasing is a preprocessor guard. Do not pass it to API calls.
const nv_dedicated_allocation_image_aliasing = 1
pub const nv_dedicated_allocation_image_aliasing_spec_version = 1
pub const nv_dedicated_allocation_image_aliasing_extension_name = "VK_NV_dedicated_allocation_image_aliasing"
// PhysicalDeviceDedicatedAllocationImageAliasingFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDedicatedAllocationImageAliasingFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    dedicated_allocation_image_aliasing Bool32
} 



// VK_EXT_buffer_device_address is a preprocessor guard. Do not pass it to API calls.
const ext_buffer_device_address = 1
pub const ext_buffer_device_address_spec_version = 2
pub const ext_buffer_device_address_extension_name = "VK_EXT_buffer_device_address"
// PhysicalDeviceBufferDeviceAddressFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceBufferDeviceAddressFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    buffer_device_address  Bool32
    buffer_device_address_capture_replay Bool32
    buffer_device_address_multi_device Bool32
} 

pub type PhysicalDeviceBufferAddressFeaturesEXT = PhysicalDeviceBufferDeviceAddressFeaturesEXT

pub type BufferDeviceAddressInfoEXT = BufferDeviceAddressInfo

// BufferDeviceAddressCreateInfoEXT extends VkBufferCreateInfo
pub struct BufferDeviceAddressCreateInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_address         DeviceAddress
} 

type VkGetBufferDeviceAddressEXT = fn (     C.Device,     &BufferDeviceAddressInfo) DeviceAddress

pub fn get_buffer_device_address_ext(
    device                                          C.Device,
    p_info                                          &BufferDeviceAddressInfo) DeviceAddress {
      f := VkGetBufferDeviceAddressEXT((*loader_p).get_sym("vkGetBufferDeviceAddressEXT"
    ) or { 
        panic("Couldn't load symbol for 'vkGetBufferDeviceAddressEXT': ${err}") })
    return f(
    device,
    p_info)
}




// VK_EXT_tooling_info is a preprocessor guard. Do not pass it to API calls.
const ext_tooling_info = 1
pub const ext_tooling_info_spec_version     = 1
pub const ext_tooling_info_extension_name   = "VK_EXT_tooling_info"
pub type ToolPurposeFlagBitsEXT = ToolPurposeFlagBits

pub type PhysicalDeviceToolPropertiesEXT = PhysicalDeviceToolProperties

type VkGetPhysicalDeviceToolPropertiesEXT = fn (     C.PhysicalDevice,     &u32,     &PhysicalDeviceToolProperties) Result

pub fn get_physical_device_tool_properties_ext(
    physical_device                                 C.PhysicalDevice,
    p_tool_count                                    &u32,
    p_tool_properties                               &PhysicalDeviceToolProperties) Result {
      f := VkGetPhysicalDeviceToolPropertiesEXT((*loader_p).get_sym('vkGetPhysicalDeviceToolPropertiesEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceToolPropertiesEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_tool_count,
    p_tool_properties)
}




// VK_EXT_separate_stencil_usage is a preprocessor guard. Do not pass it to API calls.
const ext_separate_stencil_usage = 1
pub const ext_separate_stencil_usage_spec_version = 1
pub const ext_separate_stencil_usage_extension_name = "VK_EXT_separate_stencil_usage"
pub type ImageStencilUsageCreateInfoEXT = ImageStencilUsageCreateInfo



// VK_EXT_validation_features is a preprocessor guard. Do not pass it to API calls.
const ext_validation_features = 1
pub const ext_validation_features_spec_version = 6
pub const ext_validation_features_extension_name = "VK_EXT_validation_features"

pub enum ValidationFeatureEnableEXT {
    validation_feature_enable_gpu_assisted_ext = int(0)
    validation_feature_enable_gpu_assisted_reserve_binding_slot_ext = int(1)
    validation_feature_enable_best_practices_ext = int(2)
    validation_feature_enable_debug_printf_ext = int(3)
    validation_feature_enable_synchronization_validation_ext = int(4)
    validation_feature_enable_max_enum_ext = int(0x7FFFFFFF)
}


pub enum ValidationFeatureDisableEXT {
    validation_feature_disable_all_ext = int(0)
    validation_feature_disable_shaders_ext = int(1)
    validation_feature_disable_thread_safety_ext = int(2)
    validation_feature_disable_api_parameters_ext = int(3)
    validation_feature_disable_object_lifetimes_ext = int(4)
    validation_feature_disable_core_checks_ext = int(5)
    validation_feature_disable_unique_handles_ext = int(6)
    validation_feature_disable_shader_validation_cache_ext = int(7)
    validation_feature_disable_max_enum_ext = int(0x7FFFFFFF)
}

// ValidationFeaturesEXT extends VkInstanceCreateInfo
pub struct ValidationFeaturesEXT {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    enabled_validation_feature_count            u32
    p_enabled_validation_features               &ValidationFeatureEnableEXT
    disabled_validation_feature_count           u32
    p_disabled_validation_features              &ValidationFeatureDisableEXT
} 



// VK_NV_cooperative_matrix is a preprocessor guard. Do not pass it to API calls.
const nv_cooperative_matrix = 1
pub const nv_cooperative_matrix_spec_version = 1
pub const nv_cooperative_matrix_extension_name = "VK_NV_cooperative_matrix"
pub type ComponentTypeNV = ComponentTypeKHR

pub type ScopeNV = ScopeKHR

pub struct CooperativeMatrixPropertiesNV {
mut:
    s_type                   StructureType
    p_next                   voidptr
    m_size                   u32
    n_size                   u32
    k_size                   u32
    a_type                   ComponentTypeNV
    b_type                   ComponentTypeNV
    c_type                   ComponentTypeNV
    d_type                   ComponentTypeNV
    scope                    ScopeNV
} 

// PhysicalDeviceCooperativeMatrixFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceCooperativeMatrixFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    cooperative_matrix     Bool32
    cooperative_matrix_robust_buffer_access Bool32
} 

// PhysicalDeviceCooperativeMatrixPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceCooperativeMatrixPropertiesNV {
mut:
    s_type                    StructureType
    p_next                    voidptr
    cooperative_matrix_supported_stages ShaderStageFlags
} 

type VkGetPhysicalDeviceCooperativeMatrixPropertiesNV = fn (     C.PhysicalDevice,     &u32,     &CooperativeMatrixPropertiesNV) Result

pub fn get_physical_device_cooperative_matrix_properties_nv(
    physical_device                                 C.PhysicalDevice,
    p_property_count                                &u32,
    p_properties                                    &CooperativeMatrixPropertiesNV) Result {
      f := VkGetPhysicalDeviceCooperativeMatrixPropertiesNV((*loader_p).get_sym('vkGetPhysicalDeviceCooperativeMatrixPropertiesNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceCooperativeMatrixPropertiesNV': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_property_count,
    p_properties)
}




// VK_NV_coverage_reduction_mode is a preprocessor guard. Do not pass it to API calls.
const nv_coverage_reduction_mode = 1
pub const nv_coverage_reduction_mode_spec_version = 1
pub const nv_coverage_reduction_mode_extension_name = "VK_NV_coverage_reduction_mode"

pub enum CoverageReductionModeNV {
    coverage_reduction_mode_merge_nv = int(0)
    coverage_reduction_mode_truncate_nv = int(1)
    coverage_reduction_mode_max_enum_nv = int(0x7FFFFFFF)
}

pub type PipelineCoverageReductionStateCreateFlagsNV = u32
// PhysicalDeviceCoverageReductionModeFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceCoverageReductionModeFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    coverage_reduction_mode Bool32
} 

// PipelineCoverageReductionStateCreateInfoNV extends VkPipelineMultisampleStateCreateInfo
pub struct PipelineCoverageReductionStateCreateInfoNV {
mut:
    s_type                                               StructureType
    p_next                                               voidptr
    flags                                                PipelineCoverageReductionStateCreateFlagsNV
    coverage_reduction_mode                              CoverageReductionModeNV
} 

pub struct FramebufferMixedSamplesCombinationNV {
mut:
    s_type                           StructureType
    p_next                           voidptr
    coverage_reduction_mode          CoverageReductionModeNV
    rasterization_samples            SampleCountFlagBits
    depth_stencil_samples            SampleCountFlags
    color_samples                    SampleCountFlags
} 

type VkGetPhysicalDeviceSupportedFramebufferMixedSamplesCombinationsNV = fn (     C.PhysicalDevice,     &u32,     &FramebufferMixedSamplesCombinationNV) Result

pub fn get_physical_device_supported_framebuffer_mixed_samples_combinations_nv(
    physical_device                                 C.PhysicalDevice,
    p_combination_count                             &u32,
    p_combinations                                  &FramebufferMixedSamplesCombinationNV) Result {
      f := VkGetPhysicalDeviceSupportedFramebufferMixedSamplesCombinationsNV((*loader_p).get_sym('vkGetPhysicalDeviceSupportedFramebufferMixedSamplesCombinationsNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSupportedFramebufferMixedSamplesCombinationsNV': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_combination_count,
    p_combinations)
}




// VK_EXT_fragment_shader_interlock is a preprocessor guard. Do not pass it to API calls.
const ext_fragment_shader_interlock = 1
pub const ext_fragment_shader_interlock_spec_version = 1
pub const ext_fragment_shader_interlock_extension_name = "VK_EXT_fragment_shader_interlock"
// PhysicalDeviceFragmentShaderInterlockFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceFragmentShaderInterlockFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    fragment_shader_sample_interlock Bool32
    fragment_shader_pixel_interlock Bool32
    fragment_shader_shading_rate_interlock Bool32
} 



// VK_EXT_ycbcr_image_arrays is a preprocessor guard. Do not pass it to API calls.
const ext_ycbcr_image_arrays = 1
pub const ext_ycbcr_image_arrays_spec_version = 1
pub const ext_ycbcr_image_arrays_extension_name = "VK_EXT_ycbcr_image_arrays"
// PhysicalDeviceYcbcrImageArraysFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceYcbcrImageArraysFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    ycbcr_image_arrays     Bool32
} 



// VK_EXT_provoking_vertex is a preprocessor guard. Do not pass it to API calls.
const ext_provoking_vertex = 1
pub const ext_provoking_vertex_spec_version = 1
pub const ext_provoking_vertex_extension_name = "VK_EXT_provoking_vertex"

pub enum ProvokingVertexModeEXT {
    provoking_vertex_mode_first_vertex_ext = int(0)
    provoking_vertex_mode_last_vertex_ext = int(1)
    provoking_vertex_mode_max_enum_ext = int(0x7FFFFFFF)
}

// PhysicalDeviceProvokingVertexFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceProvokingVertexFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    provoking_vertex_last  Bool32
    transform_feedback_preserves_provoking_vertex Bool32
} 

// PhysicalDeviceProvokingVertexPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceProvokingVertexPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    provoking_vertex_mode_per_pipeline Bool32
    transform_feedback_preserves_triangle_fan_provoking_vertex Bool32
} 

// PipelineRasterizationProvokingVertexStateCreateInfoEXT extends VkPipelineRasterizationStateCreateInfo
pub struct PipelineRasterizationProvokingVertexStateCreateInfoEXT {
mut:
    s_type                          StructureType
    p_next                          voidptr
    provoking_vertex_mode           ProvokingVertexModeEXT
} 



// VK_EXT_full_screen_exclusive is a preprocessor guard. Do not pass it to API calls.
const ext_full_screen_exclusive = 1
pub const ext_full_screen_exclusive_spec_version = 4
pub const ext_full_screen_exclusive_extension_name = "VK_EXT_full_screen_exclusive"

pub enum FullScreenExclusiveEXT {
    full_screen_exclusive_default_ext = int(0)
    full_screen_exclusive_allowed_ext = int(1)
    full_screen_exclusive_disallowed_ext = int(2)
    full_screen_exclusive_application_controlled_ext = int(3)
    full_screen_exclusive_max_enum_ext = int(0x7FFFFFFF)
}

// SurfaceFullScreenExclusiveInfoEXT extends VkPhysicalDeviceSurfaceInfo2KHR,VkSwapchainCreateInfoKHR
pub struct SurfaceFullScreenExclusiveInfoEXT {
mut:
    s_type                          StructureType
    p_next                          voidptr
    full_screen_exclusive           FullScreenExclusiveEXT
} 

// SurfaceCapabilitiesFullScreenExclusiveEXT extends VkSurfaceCapabilities2KHR
pub struct SurfaceCapabilitiesFullScreenExclusiveEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    full_screen_exclusive_supported Bool32
} 

// SurfaceFullScreenExclusiveWin32InfoEXT extends VkPhysicalDeviceSurfaceInfo2KHR,VkSwapchainCreateInfoKHR
pub struct SurfaceFullScreenExclusiveWin32InfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    hmonitor               voidptr
} 

type VkGetPhysicalDeviceSurfacePresentModes2EXT = fn (     C.PhysicalDevice,     &PhysicalDeviceSurfaceInfo2KHR,     &u32,     &PresentModeKHR) Result

pub fn get_physical_device_surface_present_modes2_ext(
    physical_device                                 C.PhysicalDevice,
    p_surface_info                                  &PhysicalDeviceSurfaceInfo2KHR,
    p_present_mode_count                            &u32,
    p_present_modes                                 &PresentModeKHR) Result {
      f := VkGetPhysicalDeviceSurfacePresentModes2EXT((*loader_p).get_sym('vkGetPhysicalDeviceSurfacePresentModes2EXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceSurfacePresentModes2EXT': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_surface_info,
    p_present_mode_count,
    p_present_modes)
}


type VkAcquireFullScreenExclusiveModeEXT = fn (     C.Device,     C.SwapchainKHR) Result

pub fn acquire_full_screen_exclusive_mode_ext(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR) Result {
      f := VkAcquireFullScreenExclusiveModeEXT((*loader_p).get_sym('vkAcquireFullScreenExclusiveModeEXT'
    ) or { 
        println("Couldn't load symbol for 'vkAcquireFullScreenExclusiveModeEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain)
}


type VkReleaseFullScreenExclusiveModeEXT = fn (     C.Device,     C.SwapchainKHR) Result

pub fn release_full_screen_exclusive_mode_ext(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR) Result {
      f := VkReleaseFullScreenExclusiveModeEXT((*loader_p).get_sym('vkReleaseFullScreenExclusiveModeEXT'
    ) or { 
        println("Couldn't load symbol for 'vkReleaseFullScreenExclusiveModeEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain)
}


type VkGetDeviceGroupSurfacePresentModes2EXT = fn (     C.Device,     &PhysicalDeviceSurfaceInfo2KHR,     &DeviceGroupPresentModeFlagsKHR) Result

pub fn get_device_group_surface_present_modes2_ext(
    device                                          C.Device,
    p_surface_info                                  &PhysicalDeviceSurfaceInfo2KHR,
    p_modes                                         &DeviceGroupPresentModeFlagsKHR) Result {
      f := VkGetDeviceGroupSurfacePresentModes2EXT((*loader_p).get_sym('vkGetDeviceGroupSurfacePresentModes2EXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceGroupSurfacePresentModes2EXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_surface_info,
    p_modes)
}




// VK_EXT_headless_surface is a preprocessor guard. Do not pass it to API calls.
const ext_headless_surface = 1
pub const ext_headless_surface_spec_version = 1
pub const ext_headless_surface_extension_name = "VK_EXT_headless_surface"
pub type HeadlessSurfaceCreateFlagsEXT = u32
pub struct HeadlessSurfaceCreateInfoEXT {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    flags                                  HeadlessSurfaceCreateFlagsEXT
} 

type VkCreateHeadlessSurfaceEXT = fn (     C.Instance,     &HeadlessSurfaceCreateInfoEXT,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_headless_surface_ext(
    instance                                        C.Instance,
    p_create_info                                   &HeadlessSurfaceCreateInfoEXT,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateHeadlessSurfaceEXT((*loader_p).get_sym('vkCreateHeadlessSurfaceEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCreateHeadlessSurfaceEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}




// VK_EXT_line_rasterization is a preprocessor guard. Do not pass it to API calls.
const ext_line_rasterization = 1
pub const ext_line_rasterization_spec_version = 1
pub const ext_line_rasterization_extension_name = "VK_EXT_line_rasterization"

pub enum LineRasterizationModeEXT {
    line_rasterization_mode_default_ext = int(0)
    line_rasterization_mode_rectangular_ext = int(1)
    line_rasterization_mode_bresenham_ext = int(2)
    line_rasterization_mode_rectangular_smooth_ext = int(3)
    line_rasterization_mode_max_enum_ext = int(0x7FFFFFFF)
}

// PhysicalDeviceLineRasterizationFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceLineRasterizationFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    rectangular_lines      Bool32
    bresenham_lines        Bool32
    smooth_lines           Bool32
    stippled_rectangular_lines Bool32
    stippled_bresenham_lines Bool32
    stippled_smooth_lines  Bool32
} 

// PhysicalDeviceLineRasterizationPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceLineRasterizationPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    line_sub_pixel_precision_bits u32
} 

// PipelineRasterizationLineStateCreateInfoEXT extends VkPipelineRasterizationStateCreateInfo
pub struct PipelineRasterizationLineStateCreateInfoEXT {
mut:
    s_type                            StructureType
    p_next                            voidptr
    line_rasterization_mode           LineRasterizationModeEXT
    stippled_line_enable              Bool32
    line_stipple_factor               u32
    line_stipple_pattern              u16
} 

type VkCmdSetLineStippleEXT = fn (     C.CommandBuffer,     u32,     u16) 

pub fn cmd_set_line_stipple_ext(
    command_buffer                                  C.CommandBuffer,
    line_stipple_factor                             u32,
    line_stipple_pattern                            u16)  {
      f := VkCmdSetLineStippleEXT((*loader_p).get_sym('vkCmdSetLineStippleEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetLineStippleEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    line_stipple_factor,
    line_stipple_pattern)
}




// VK_EXT_shader_atomic_float is a preprocessor guard. Do not pass it to API calls.
const ext_shader_atomic_float = 1
pub const ext_shader_atomic_float_spec_version = 1
pub const ext_shader_atomic_float_extension_name = "VK_EXT_shader_atomic_float"
// PhysicalDeviceShaderAtomicFloatFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderAtomicFloatFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_buffer_float32_atomics Bool32
    shader_buffer_float32_atomic_add Bool32
    shader_buffer_float64_atomics Bool32
    shader_buffer_float64_atomic_add Bool32
    shader_shared_float32_atomics Bool32
    shader_shared_float32_atomic_add Bool32
    shader_shared_float64_atomics Bool32
    shader_shared_float64_atomic_add Bool32
    shader_image_float32_atomics Bool32
    shader_image_float32_atomic_add Bool32
    sparse_image_float32_atomics Bool32
    sparse_image_float32_atomic_add Bool32
} 



// VK_EXT_host_query_reset is a preprocessor guard. Do not pass it to API calls.
const ext_host_query_reset = 1
pub const ext_host_query_reset_spec_version = 1
pub const ext_host_query_reset_extension_name = "VK_EXT_host_query_reset"
pub type PhysicalDeviceHostQueryResetFeaturesEXT = PhysicalDeviceHostQueryResetFeatures

type VkResetQueryPoolEXT = fn (     C.Device,     C.QueryPool,     u32,     u32) 

pub fn reset_query_pool_ext(
    device                                          C.Device,
    query_pool                                      C.QueryPool,
    first_query                                     u32,
    query_count                                     u32)  {
      f := VkResetQueryPoolEXT((*loader_p).get_sym('vkResetQueryPoolEXT'
    ) or { 
        println("Couldn't load symbol for 'vkResetQueryPoolEXT': ${err}")
        return 
    })
    f(
    device,
    query_pool,
    first_query,
    query_count)
}




// VK_EXT_index_type_uint8 is a preprocessor guard. Do not pass it to API calls.
const ext_index_type_uint8 = 1
pub const ext_index_type_uint8_spec_version = 1
pub const ext_index_type_uint8_extension_name = "VK_EXT_index_type_uint8"
// PhysicalDeviceIndexTypeUint8FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceIndexTypeUint8FeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    index_type_uint8       Bool32
} 



// VK_EXT_extended_dynamic_state is a preprocessor guard. Do not pass it to API calls.
const ext_extended_dynamic_state = 1
pub const ext_extended_dynamic_state_spec_version = 1
pub const ext_extended_dynamic_state_extension_name = "VK_EXT_extended_dynamic_state"
// PhysicalDeviceExtendedDynamicStateFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceExtendedDynamicStateFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    extended_dynamic_state Bool32
} 

type VkCmdSetCullModeEXT = fn (     C.CommandBuffer,     CullModeFlags) 

pub fn cmd_set_cull_mode_ext(
    command_buffer                                  C.CommandBuffer,
    cull_mode                                       CullModeFlags)  {
      f := VkCmdSetCullModeEXT((*loader_p).get_sym('vkCmdSetCullModeEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetCullModeEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    cull_mode)
}


type VkCmdSetFrontFaceEXT = fn (     C.CommandBuffer,     FrontFace) 

pub fn cmd_set_front_face_ext(
    command_buffer                                  C.CommandBuffer,
    front_face                                      FrontFace)  {
      f := VkCmdSetFrontFaceEXT((*loader_p).get_sym('vkCmdSetFrontFaceEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetFrontFaceEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    front_face)
}


type VkCmdSetPrimitiveTopologyEXT = fn (     C.CommandBuffer,     PrimitiveTopology) 

pub fn cmd_set_primitive_topology_ext(
    command_buffer                                  C.CommandBuffer,
    primitive_topology                              PrimitiveTopology)  {
      f := VkCmdSetPrimitiveTopologyEXT((*loader_p).get_sym('vkCmdSetPrimitiveTopologyEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetPrimitiveTopologyEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    primitive_topology)
}


type VkCmdSetViewportWithCountEXT = fn (     C.CommandBuffer,     u32,     &Viewport) 

pub fn cmd_set_viewport_with_count_ext(
    command_buffer                                  C.CommandBuffer,
    viewport_count                                  u32,
    p_viewports                                     &Viewport)  {
      f := VkCmdSetViewportWithCountEXT((*loader_p).get_sym('vkCmdSetViewportWithCountEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetViewportWithCountEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    viewport_count,
    p_viewports)
}


type VkCmdSetScissorWithCountEXT = fn (     C.CommandBuffer,     u32,     &Rect2D) 

pub fn cmd_set_scissor_with_count_ext(
    command_buffer                                  C.CommandBuffer,
    scissor_count                                   u32,
    p_scissors                                      &Rect2D)  {
      f := VkCmdSetScissorWithCountEXT((*loader_p).get_sym('vkCmdSetScissorWithCountEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetScissorWithCountEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    scissor_count,
    p_scissors)
}


type VkCmdBindVertexBuffers2EXT = fn (     C.CommandBuffer,     u32,     u32,     &C.Buffer,     &DeviceSize,     &DeviceSize,     &DeviceSize) 

pub fn cmd_bind_vertex_buffers2_ext(
    command_buffer                                  C.CommandBuffer,
    first_binding                                   u32,
    binding_count                                   u32,
    p_buffers                                       &C.Buffer,
    p_offsets                                       &DeviceSize,
    p_sizes                                         &DeviceSize,
    p_strides                                       &DeviceSize)  {
      f := VkCmdBindVertexBuffers2EXT((*loader_p).get_sym('vkCmdBindVertexBuffers2EXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindVertexBuffers2EXT': ${err}")
        return 
    })
    f(
    command_buffer,
    first_binding,
    binding_count,
    p_buffers,
    p_offsets,
    p_sizes,
    p_strides)
}


type VkCmdSetDepthTestEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_depth_test_enable_ext(
    command_buffer                                  C.CommandBuffer,
    depth_test_enable                               Bool32)  {
      f := VkCmdSetDepthTestEnableEXT((*loader_p).get_sym('vkCmdSetDepthTestEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthTestEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_test_enable)
}


type VkCmdSetDepthWriteEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_depth_write_enable_ext(
    command_buffer                                  C.CommandBuffer,
    depth_write_enable                              Bool32)  {
      f := VkCmdSetDepthWriteEnableEXT((*loader_p).get_sym('vkCmdSetDepthWriteEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthWriteEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_write_enable)
}


type VkCmdSetDepthCompareOpEXT = fn (     C.CommandBuffer,     CompareOp) 

pub fn cmd_set_depth_compare_op_ext(
    command_buffer                                  C.CommandBuffer,
    depth_compare_op                                CompareOp)  {
      f := VkCmdSetDepthCompareOpEXT((*loader_p).get_sym('vkCmdSetDepthCompareOpEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthCompareOpEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_compare_op)
}


type VkCmdSetDepthBoundsTestEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_depth_bounds_test_enable_ext(
    command_buffer                                  C.CommandBuffer,
    depth_bounds_test_enable                        Bool32)  {
      f := VkCmdSetDepthBoundsTestEnableEXT((*loader_p).get_sym('vkCmdSetDepthBoundsTestEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthBoundsTestEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_bounds_test_enable)
}


type VkCmdSetStencilTestEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_stencil_test_enable_ext(
    command_buffer                                  C.CommandBuffer,
    stencil_test_enable                             Bool32)  {
      f := VkCmdSetStencilTestEnableEXT((*loader_p).get_sym('vkCmdSetStencilTestEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetStencilTestEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    stencil_test_enable)
}


type VkCmdSetStencilOpEXT = fn (     C.CommandBuffer,     StencilFaceFlags,     StencilOp,     StencilOp,     StencilOp,     CompareOp) 

pub fn cmd_set_stencil_op_ext(
    command_buffer                                  C.CommandBuffer,
    face_mask                                       StencilFaceFlags,
    fail_op                                         StencilOp,
    pass_op                                         StencilOp,
    depth_fail_op                                   StencilOp,
    compare_op                                      CompareOp)  {
      f := VkCmdSetStencilOpEXT((*loader_p).get_sym('vkCmdSetStencilOpEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetStencilOpEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    face_mask,
    fail_op,
    pass_op,
    depth_fail_op,
    compare_op)
}




// VK_EXT_host_image_copy is a preprocessor guard. Do not pass it to API calls.
const ext_host_image_copy = 1
pub const ext_host_image_copy_spec_version  = 1
pub const ext_host_image_copy_extension_name = "VK_EXT_host_image_copy"

pub enum HostImageCopyFlagBitsEXT {
    host_image_copy_memcpy_ext = int(0x00000001)
    host_image_copy_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type HostImageCopyFlagsEXT = u32
// PhysicalDeviceHostImageCopyFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceHostImageCopyFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    host_image_copy        Bool32
} 

// PhysicalDeviceHostImageCopyPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceHostImageCopyPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    copy_src_layout_count  u32
    p_copy_src_layouts     &ImageLayout
    copy_dst_layout_count  u32
    p_copy_dst_layouts     &ImageLayout
    optimal_tiling_layout_uuid []u8
    identical_memory_type_requirements Bool32
} 

pub struct MemoryToImageCopyEXT {
mut:
    s_type                          StructureType
    p_next                          voidptr
    p_host_pointer                  voidptr
    memory_row_length               u32
    memory_image_height             u32
    image_subresource               ImageSubresourceLayers
    image_offset                    Offset3D
    image_extent                    Extent3D
} 

pub struct ImageToMemoryCopyEXT {
mut:
    s_type                          StructureType
    p_next                          voidptr
    p_host_pointer                  voidptr
    memory_row_length               u32
    memory_image_height             u32
    image_subresource               ImageSubresourceLayers
    image_offset                    Offset3D
    image_extent                    Extent3D
} 

pub struct CopyMemoryToImageInfoEXT {
mut:
    s_type                               StructureType
    p_next                               voidptr
    flags                                HostImageCopyFlagsEXT
    dst_image                            C.Image
    dst_image_layout                     ImageLayout
    region_count                         u32
    p_regions                            &MemoryToImageCopyEXT
} 

pub struct CopyImageToMemoryInfoEXT {
mut:
    s_type                               StructureType
    p_next                               voidptr
    flags                                HostImageCopyFlagsEXT
    src_image                            C.Image
    src_image_layout                     ImageLayout
    region_count                         u32
    p_regions                            &ImageToMemoryCopyEXT
} 

pub struct CopyImageToImageInfoEXT {
mut:
    s_type                         StructureType
    p_next                         voidptr
    flags                          HostImageCopyFlagsEXT
    src_image                      C.Image
    src_image_layout               ImageLayout
    dst_image                      C.Image
    dst_image_layout               ImageLayout
    region_count                   u32
    p_regions                      &ImageCopy2
} 

pub struct HostImageLayoutTransitionInfoEXT {
mut:
    s_type                         StructureType
    p_next                         voidptr
    image                          C.Image
    old_layout                     ImageLayout
    new_layout                     ImageLayout
    subresource_range              ImageSubresourceRange
} 

// SubresourceHostMemcpySizeEXT extends VkSubresourceLayout2KHR
pub struct SubresourceHostMemcpySizeEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    size                   DeviceSize
} 

// HostImageCopyDevicePerformanceQueryEXT extends VkImageFormatProperties2
pub struct HostImageCopyDevicePerformanceQueryEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    optimal_device_access  Bool32
    identical_memory_layout Bool32
} 

pub type SubresourceLayout2EXT = SubresourceLayout2KHR

pub type ImageSubresource2EXT = ImageSubresource2KHR

type VkCopyMemoryToImageEXT = fn (     C.Device,     &CopyMemoryToImageInfoEXT) Result

pub fn copy_memory_to_image_ext(
    device                                          C.Device,
    p_copy_memory_to_image_info                     &CopyMemoryToImageInfoEXT) Result {
      f := VkCopyMemoryToImageEXT((*loader_p).get_sym('vkCopyMemoryToImageEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCopyMemoryToImageEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_copy_memory_to_image_info)
}


type VkCopyImageToMemoryEXT = fn (     C.Device,     &CopyImageToMemoryInfoEXT) Result

pub fn copy_image_to_memory_ext(
    device                                          C.Device,
    p_copy_image_to_memory_info                     &CopyImageToMemoryInfoEXT) Result {
      f := VkCopyImageToMemoryEXT((*loader_p).get_sym('vkCopyImageToMemoryEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCopyImageToMemoryEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_copy_image_to_memory_info)
}


type VkCopyImageToImageEXT = fn (     C.Device,     &CopyImageToImageInfoEXT) Result

pub fn copy_image_to_image_ext(
    device                                          C.Device,
    p_copy_image_to_image_info                      &CopyImageToImageInfoEXT) Result {
      f := VkCopyImageToImageEXT((*loader_p).get_sym('vkCopyImageToImageEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCopyImageToImageEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_copy_image_to_image_info)
}


type VkTransitionImageLayoutEXT = fn (     C.Device,     u32,     &HostImageLayoutTransitionInfoEXT) Result

pub fn transition_image_layout_ext(
    device                                          C.Device,
    transition_count                                u32,
    p_transitions                                   &HostImageLayoutTransitionInfoEXT) Result {
      f := VkTransitionImageLayoutEXT((*loader_p).get_sym('vkTransitionImageLayoutEXT'
    ) or { 
        println("Couldn't load symbol for 'vkTransitionImageLayoutEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    transition_count,
    p_transitions)
}


type VkGetImageSubresourceLayout2EXT = fn (     C.Device,     C.Image,     &ImageSubresource2KHR,     &SubresourceLayout2KHR) 

pub fn get_image_subresource_layout2_ext(
    device                                          C.Device,
    image                                           C.Image,
    p_subresource                                   &ImageSubresource2KHR,
    p_layout                                        &SubresourceLayout2KHR)  {
      f := VkGetImageSubresourceLayout2EXT((*loader_p).get_sym('vkGetImageSubresourceLayout2EXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageSubresourceLayout2EXT': ${err}")
        return 
    })
    f(
    device,
    image,
    p_subresource,
    p_layout)
}




// VK_EXT_shader_atomic_float2 is a preprocessor guard. Do not pass it to API calls.
const ext_shader_atomic_float2 = 1
pub const ext_shader_atomic_float_2_spec_version = 1
pub const ext_shader_atomic_float_2_extension_name = "VK_EXT_shader_atomic_float2"
// PhysicalDeviceShaderAtomicFloat2FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderAtomicFloat2FeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_buffer_float16_atomics Bool32
    shader_buffer_float16_atomic_add Bool32
    shader_buffer_float16_atomic_min_max Bool32
    shader_buffer_float32_atomic_min_max Bool32
    shader_buffer_float64_atomic_min_max Bool32
    shader_shared_float16_atomics Bool32
    shader_shared_float16_atomic_add Bool32
    shader_shared_float16_atomic_min_max Bool32
    shader_shared_float32_atomic_min_max Bool32
    shader_shared_float64_atomic_min_max Bool32
    shader_image_float32_atomic_min_max Bool32
    sparse_image_float32_atomic_min_max Bool32
} 



// VK_EXT_surface_maintenance1 is a preprocessor guard. Do not pass it to API calls.
const ext_surface_maintenance1 = 1
pub const ext_surface_maintenance_1_spec_version = 1
pub const ext_surface_maintenance_1_extension_name = "VK_EXT_surface_maintenance1"

pub enum PresentScalingFlagBitsEXT {
    present_scaling_one_to_one_bit_ext = int(0x00000001)
    present_scaling_aspect_ratio_stretch_bit_ext = int(0x00000002)
    present_scaling_stretch_bit_ext = int(0x00000004)
    present_scaling_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type PresentScalingFlagsEXT = u32

pub enum PresentGravityFlagBitsEXT {
    present_gravity_min_bit_ext = int(0x00000001)
    present_gravity_max_bit_ext = int(0x00000002)
    present_gravity_centered_bit_ext = int(0x00000004)
    present_gravity_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type PresentGravityFlagsEXT = u32
// SurfacePresentModeEXT extends VkPhysicalDeviceSurfaceInfo2KHR
pub struct SurfacePresentModeEXT {
mut:
    s_type                  StructureType
    p_next                  voidptr
    present_mode            PresentModeKHR
} 

// SurfacePresentScalingCapabilitiesEXT extends VkSurfaceCapabilities2KHR
pub struct SurfacePresentScalingCapabilitiesEXT {
mut:
    s_type                          StructureType
    p_next                          voidptr
    supported_present_scaling       PresentScalingFlagsEXT
    supported_present_gravity_x     PresentGravityFlagsEXT
    supported_present_gravity_y     PresentGravityFlagsEXT
    min_scaled_image_extent         Extent2D
    max_scaled_image_extent         Extent2D
} 

// SurfacePresentModeCompatibilityEXT extends VkSurfaceCapabilities2KHR
pub struct SurfacePresentModeCompatibilityEXT {
mut:
    s_type                   StructureType
    p_next                   voidptr
    present_mode_count       u32
    p_present_modes          &PresentModeKHR
} 



// VK_EXT_swapchain_maintenance1 is a preprocessor guard. Do not pass it to API calls.
const ext_swapchain_maintenance1 = 1
pub const ext_swapchain_maintenance_1_spec_version = 1
pub const ext_swapchain_maintenance_1_extension_name = "VK_EXT_swapchain_maintenance1"
// PhysicalDeviceSwapchainMaintenance1FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceSwapchainMaintenance1FeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    swapchain_maintenance1 Bool32
} 

// SwapchainPresentFenceInfoEXT extends VkPresentInfoKHR
pub struct SwapchainPresentFenceInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    swapchain_count        u32
    p_fences               &C.Fence
} 

// SwapchainPresentModesCreateInfoEXT extends VkSwapchainCreateInfoKHR
pub struct SwapchainPresentModesCreateInfoEXT {
mut:
    s_type                         StructureType
    p_next                         voidptr
    present_mode_count             u32
    p_present_modes                &PresentModeKHR
} 

// SwapchainPresentModeInfoEXT extends VkPresentInfoKHR
pub struct SwapchainPresentModeInfoEXT {
mut:
    s_type                         StructureType
    p_next                         voidptr
    swapchain_count                u32
    p_present_modes                &PresentModeKHR
} 

// SwapchainPresentScalingCreateInfoEXT extends VkSwapchainCreateInfoKHR
pub struct SwapchainPresentScalingCreateInfoEXT {
mut:
    s_type                          StructureType
    p_next                          voidptr
    scaling_behavior                PresentScalingFlagsEXT
    present_gravity_x               PresentGravityFlagsEXT
    present_gravity_y               PresentGravityFlagsEXT
} 

pub struct ReleaseSwapchainImagesInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    swapchain              C.SwapchainKHR
    image_index_count      u32
    p_image_indices        &u32
} 

type VkReleaseSwapchainImagesEXT = fn (     C.Device,     &ReleaseSwapchainImagesInfoEXT) Result

pub fn release_swapchain_images_ext(
    device                                          C.Device,
    p_release_info                                  &ReleaseSwapchainImagesInfoEXT) Result {
      f := VkReleaseSwapchainImagesEXT((*loader_p).get_sym('vkReleaseSwapchainImagesEXT'
    ) or { 
        println("Couldn't load symbol for 'vkReleaseSwapchainImagesEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_release_info)
}




// VK_EXT_shader_demote_to_helper_invocation is a preprocessor guard. Do not pass it to API calls.
const ext_shader_demote_to_helper_invocation = 1
pub const ext_shader_demote_to_helper_invocation_spec_version = 1
pub const ext_shader_demote_to_helper_invocation_extension_name = "VK_EXT_shader_demote_to_helper_invocation"
pub type PhysicalDeviceShaderDemoteToHelperInvocationFeaturesEXT = PhysicalDeviceShaderDemoteToHelperInvocationFeatures



// VK_NV_device_generated_commands is a preprocessor guard. Do not pass it to API calls.
const nv_device_generated_commands = 1
pub type C.IndirectCommandsLayoutNV = voidptr
pub const nv_device_generated_commands_spec_version = 3
pub const nv_device_generated_commands_extension_name = "VK_NV_device_generated_commands"

pub enum IndirectCommandsTokenTypeNV {
    indirect_commands_token_type_shader_group_nv = int(0)
    indirect_commands_token_type_state_flags_nv = int(1)
    indirect_commands_token_type_index_buffer_nv = int(2)
    indirect_commands_token_type_vertex_buffer_nv = int(3)
    indirect_commands_token_type_push_constant_nv = int(4)
    indirect_commands_token_type_draw_indexed_nv = int(5)
    indirect_commands_token_type_draw_nv = int(6)
    indirect_commands_token_type_draw_tasks_nv = int(7)
    indirect_commands_token_type_draw_mesh_tasks_nv = int(1000328000)
    indirect_commands_token_type_pipeline_nv = int(1000428003)
    indirect_commands_token_type_dispatch_nv = int(1000428004)
    indirect_commands_token_type_max_enum_nv = int(0x7FFFFFFF)
}


pub enum IndirectStateFlagBitsNV {
    indirect_state_flag_frontface_bit_nv = int(0x00000001)
    indirect_state_flag_bits_max_enum_nv = int(0x7FFFFFFF)
}

pub type IndirectStateFlagsNV = u32

pub enum IndirectCommandsLayoutUsageFlagBitsNV {
    indirect_commands_layout_usage_explicit_preprocess_bit_nv = int(0x00000001)
    indirect_commands_layout_usage_indexed_sequences_bit_nv = int(0x00000002)
    indirect_commands_layout_usage_unordered_sequences_bit_nv = int(0x00000004)
    indirect_commands_layout_usage_flag_bits_max_enum_nv = int(0x7FFFFFFF)
}

pub type IndirectCommandsLayoutUsageFlagsNV = u32
// PhysicalDeviceDeviceGeneratedCommandsPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceDeviceGeneratedCommandsPropertiesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_graphics_shader_group_count u32
    max_indirect_sequence_count u32
    max_indirect_commands_token_count u32
    max_indirect_commands_stream_count u32
    max_indirect_commands_token_offset u32
    max_indirect_commands_stream_stride u32
    min_sequences_count_buffer_offset_alignment u32
    min_sequences_index_buffer_offset_alignment u32
    min_indirect_commands_buffer_offset_alignment u32
} 

// PhysicalDeviceDeviceGeneratedCommandsFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDeviceGeneratedCommandsFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_generated_commands Bool32
} 

pub struct GraphicsShaderGroupCreateInfoNV {
mut:
    s_type                                              StructureType
    p_next                                              voidptr
    stage_count                                         u32
    p_stages                                            &PipelineShaderStageCreateInfo
    p_vertex_input_state                                &PipelineVertexInputStateCreateInfo
    p_tessellation_state                                &PipelineTessellationStateCreateInfo
} 

// GraphicsPipelineShaderGroupsCreateInfoNV extends VkGraphicsPipelineCreateInfo
pub struct GraphicsPipelineShaderGroupsCreateInfoNV {
mut:
    s_type                                          StructureType
    p_next                                          voidptr
    group_count                                     u32
    p_groups                                        &GraphicsShaderGroupCreateInfoNV
    pipeline_count                                  u32
    p_pipelines                                     &C.Pipeline
} 

pub struct BindShaderGroupIndirectCommandNV {
mut:
    group_index     u32
} 

pub struct BindIndexBufferIndirectCommandNV {
mut:
    buffer_address         DeviceAddress
    size                   u32
    index_type             IndexType
} 

pub struct BindVertexBufferIndirectCommandNV {
mut:
    buffer_address         DeviceAddress
    size                   u32
    stride                 u32
} 

pub struct SetStateFlagsIndirectCommandNV {
mut:
    data            u32
} 

pub struct IndirectCommandsStreamNV {
mut:
    buffer              C.Buffer
    offset              DeviceSize
} 

pub struct IndirectCommandsLayoutTokenNV {
mut:
    s_type                               StructureType
    p_next                               voidptr
    token_type                           IndirectCommandsTokenTypeNV
    stream                               u32
    offset                               u32
    vertex_binding_unit                  u32
    vertex_dynamic_stride                Bool32
    pushconstant_pipeline_layout         C.PipelineLayout
    pushconstant_shader_stage_flags      ShaderStageFlags
    pushconstant_offset                  u32
    pushconstant_size                    u32
    indirect_state_flags                 IndirectStateFlagsNV
    index_type_count                     u32
    p_index_types                        &IndexType
    p_index_type_values                  &u32
} 

pub struct IndirectCommandsLayoutCreateInfoNV {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    flags                                         IndirectCommandsLayoutUsageFlagsNV
    pipeline_bind_point                           PipelineBindPoint
    token_count                                   u32
    p_tokens                                      &IndirectCommandsLayoutTokenNV
    stream_count                                  u32
    p_stream_strides                              &u32
} 

pub struct GeneratedCommandsInfoNV {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    pipeline_bind_point                      PipelineBindPoint
    pipeline                                 C.Pipeline
    indirect_commands_layout                 C.IndirectCommandsLayoutNV
    stream_count                             u32
    p_streams                                &IndirectCommandsStreamNV
    sequences_count                          u32
    preprocess_buffer                        C.Buffer
    preprocess_offset                        DeviceSize
    preprocess_size                          DeviceSize
    sequences_count_buffer                   C.Buffer
    sequences_count_offset                   DeviceSize
    sequences_index_buffer                   C.Buffer
    sequences_index_offset                   DeviceSize
} 

pub struct GeneratedCommandsMemoryRequirementsInfoNV {
mut:
    s_type                            StructureType
    p_next                            voidptr
    pipeline_bind_point               PipelineBindPoint
    pipeline                          C.Pipeline
    indirect_commands_layout          C.IndirectCommandsLayoutNV
    max_sequences_count               u32
} 

type VkGetGeneratedCommandsMemoryRequirementsNV = fn (     C.Device,     &GeneratedCommandsMemoryRequirementsInfoNV,     &MemoryRequirements2) 

pub fn get_generated_commands_memory_requirements_nv(
    device                                          C.Device,
    p_info                                          &GeneratedCommandsMemoryRequirementsInfoNV,
    p_memory_requirements                           &MemoryRequirements2)  {
      f := VkGetGeneratedCommandsMemoryRequirementsNV((*loader_p).get_sym('vkGetGeneratedCommandsMemoryRequirementsNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetGeneratedCommandsMemoryRequirementsNV': ${err}")
        return 
    })
    f(
    device,
    p_info,
    p_memory_requirements)
}


type VkCmdPreprocessGeneratedCommandsNV = fn (     C.CommandBuffer,     &GeneratedCommandsInfoNV) 

pub fn cmd_preprocess_generated_commands_nv(
    command_buffer                                  C.CommandBuffer,
    p_generated_commands_info                       &GeneratedCommandsInfoNV)  {
      f := VkCmdPreprocessGeneratedCommandsNV((*loader_p).get_sym('vkCmdPreprocessGeneratedCommandsNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdPreprocessGeneratedCommandsNV': ${err}")
        return 
    })
    f(
    command_buffer,
    p_generated_commands_info)
}


type VkCmdExecuteGeneratedCommandsNV = fn (     C.CommandBuffer,     Bool32,     &GeneratedCommandsInfoNV) 

pub fn cmd_execute_generated_commands_nv(
    command_buffer                                  C.CommandBuffer,
    is_preprocessed                                 Bool32,
    p_generated_commands_info                       &GeneratedCommandsInfoNV)  {
      f := VkCmdExecuteGeneratedCommandsNV((*loader_p).get_sym('vkCmdExecuteGeneratedCommandsNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdExecuteGeneratedCommandsNV': ${err}")
        return 
    })
    f(
    command_buffer,
    is_preprocessed,
    p_generated_commands_info)
}


type VkCmdBindPipelineShaderGroupNV = fn (     C.CommandBuffer,     PipelineBindPoint,     C.Pipeline,     u32) 

pub fn cmd_bind_pipeline_shader_group_nv(
    command_buffer                                  C.CommandBuffer,
    pipeline_bind_point                             PipelineBindPoint,
    pipeline                                        C.Pipeline,
    group_index                                     u32)  {
      f := VkCmdBindPipelineShaderGroupNV((*loader_p).get_sym('vkCmdBindPipelineShaderGroupNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindPipelineShaderGroupNV': ${err}")
        return 
    })
    f(
    command_buffer,
    pipeline_bind_point,
    pipeline,
    group_index)
}


type VkCreateIndirectCommandsLayoutNV = fn (     C.Device,     &IndirectCommandsLayoutCreateInfoNV,     &AllocationCallbacks,     &C.IndirectCommandsLayoutNV) Result

pub fn create_indirect_commands_layout_nv(
    device                                          C.Device,
    p_create_info                                   &IndirectCommandsLayoutCreateInfoNV,
    p_allocator                                     &AllocationCallbacks,
    p_indirect_commands_layout                      &C.IndirectCommandsLayoutNV) Result {
      f := VkCreateIndirectCommandsLayoutNV((*loader_p).get_sym('vkCreateIndirectCommandsLayoutNV'
    ) or { 
        println("Couldn't load symbol for 'vkCreateIndirectCommandsLayoutNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_indirect_commands_layout)
}


type VkDestroyIndirectCommandsLayoutNV = fn (     C.Device,     C.IndirectCommandsLayoutNV,     &AllocationCallbacks) 

pub fn destroy_indirect_commands_layout_nv(
    device                                          C.Device,
    indirect_commands_layout                        C.IndirectCommandsLayoutNV,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyIndirectCommandsLayoutNV((*loader_p).get_sym('vkDestroyIndirectCommandsLayoutNV'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyIndirectCommandsLayoutNV': ${err}")
        return 
    })
    f(
    device,
    indirect_commands_layout,
    p_allocator)
}




// VK_NV_inherited_viewport_scissor is a preprocessor guard. Do not pass it to API calls.
const nv_inherited_viewport_scissor = 1
pub const nv_inherited_viewport_scissor_spec_version = 1
pub const nv_inherited_viewport_scissor_extension_name = "VK_NV_inherited_viewport_scissor"
// PhysicalDeviceInheritedViewportScissorFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceInheritedViewportScissorFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    inherited_viewport_scissor2_d Bool32
} 

// CommandBufferInheritanceViewportScissorInfoNV extends VkCommandBufferInheritanceInfo
pub struct CommandBufferInheritanceViewportScissorInfoNV {
mut:
    s_type                   StructureType
    p_next                   voidptr
    viewport_scissor2_d      Bool32
    viewport_depth_count     u32
    p_viewport_depths        &Viewport
} 



// VK_EXT_texel_buffer_alignment is a preprocessor guard. Do not pass it to API calls.
const ext_texel_buffer_alignment = 1
pub const ext_texel_buffer_alignment_spec_version = 1
pub const ext_texel_buffer_alignment_extension_name = "VK_EXT_texel_buffer_alignment"
// PhysicalDeviceTexelBufferAlignmentFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceTexelBufferAlignmentFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    texel_buffer_alignment Bool32
} 

pub type PhysicalDeviceTexelBufferAlignmentPropertiesEXT = PhysicalDeviceTexelBufferAlignmentProperties



// VK_QCOM_render_pass_transform is a preprocessor guard. Do not pass it to API calls.
const qcom_render_pass_transform = 1
pub const qcom_render_pass_transform_spec_version = 3
pub const qcom_render_pass_transform_extension_name = "VK_QCOM_render_pass_transform"
// RenderPassTransformBeginInfoQCOM extends VkRenderPassBeginInfo
pub struct RenderPassTransformBeginInfoQCOM {
mut:
    s_type                               StructureType
    p_next                               voidptr
    transform                            SurfaceTransformFlagBitsKHR
} 

// CommandBufferInheritanceRenderPassTransformInfoQCOM extends VkCommandBufferInheritanceInfo
pub struct CommandBufferInheritanceRenderPassTransformInfoQCOM {
mut:
    s_type                               StructureType
    p_next                               voidptr
    transform                            SurfaceTransformFlagBitsKHR
    render_area                          Rect2D
} 



// VK_EXT_depth_bias_control is a preprocessor guard. Do not pass it to API calls.
const ext_depth_bias_control = 1
pub const ext_depth_bias_control_spec_version = 1
pub const ext_depth_bias_control_extension_name = "VK_EXT_depth_bias_control"

pub enum DepthBiasRepresentationEXT {
    depth_bias_representation_least_representable_value_format_ext = int(0)
    depth_bias_representation_least_representable_value_force_unorm_ext = int(1)
    depth_bias_representation_float_ext = int(2)
    depth_bias_representation_max_enum_ext = int(0x7FFFFFFF)
}

// PhysicalDeviceDepthBiasControlFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDepthBiasControlFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    depth_bias_control     Bool32
    least_representable_value_force_unorm_representation Bool32
    float_representation   Bool32
    depth_bias_exact       Bool32
} 

pub struct DepthBiasInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    depth_bias_constant_factor f32
    depth_bias_clamp       f32
    depth_bias_slope_factor f32
} 

// DepthBiasRepresentationInfoEXT extends VkDepthBiasInfoEXT,VkPipelineRasterizationStateCreateInfo
pub struct DepthBiasRepresentationInfoEXT {
mut:
    s_type                              StructureType
    p_next                              voidptr
    depth_bias_representation           DepthBiasRepresentationEXT
    depth_bias_exact                    Bool32
} 

type VkCmdSetDepthBias2EXT = fn (     C.CommandBuffer,     &DepthBiasInfoEXT) 

pub fn cmd_set_depth_bias2_ext(
    command_buffer                                  C.CommandBuffer,
    p_depth_bias_info                               &DepthBiasInfoEXT)  {
      f := VkCmdSetDepthBias2EXT((*loader_p).get_sym('vkCmdSetDepthBias2EXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthBias2EXT': ${err}")
        return 
    })
    f(
    command_buffer,
    p_depth_bias_info)
}




// VK_EXT_device_memory_report is a preprocessor guard. Do not pass it to API calls.
const ext_device_memory_report = 1
pub const ext_device_memory_report_spec_version = 2
pub const ext_device_memory_report_extension_name = "VK_EXT_device_memory_report"

pub enum DeviceMemoryReportEventTypeEXT {
    device_memory_report_event_type_allocate_ext = int(0)
    device_memory_report_event_type_free_ext = int(1)
    device_memory_report_event_type_import_ext = int(2)
    device_memory_report_event_type_unimport_ext = int(3)
    device_memory_report_event_type_allocation_failed_ext = int(4)
    device_memory_report_event_type_max_enum_ext = int(0x7FFFFFFF)
}

pub type DeviceMemoryReportFlagsEXT = u32
// PhysicalDeviceDeviceMemoryReportFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDeviceMemoryReportFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_memory_report   Bool32
} 

pub struct DeviceMemoryReportCallbackDataEXT {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    flags                                   DeviceMemoryReportFlagsEXT
    vktype                                  DeviceMemoryReportEventTypeEXT
    memory_object_id                        u64
    size                                    DeviceSize
    object_type                             ObjectType
    object_handle                           u64
    heap_index                              u32
} 

pub type PFN_vkDeviceMemoryReportCallbackEXT = fn (   pCallbackData                     &DeviceMemoryReportCallbackDataEXT,   pUserData                         voidptr) voidptr
// DeviceDeviceMemoryReportCreateInfoEXT extends VkDeviceCreateInfo
pub struct DeviceDeviceMemoryReportCreateInfoEXT {
mut:
    s_type                                     StructureType
    p_next                                     voidptr
    flags                                      DeviceMemoryReportFlagsEXT
    pfn_user_callback                          PFN_vkDeviceMemoryReportCallbackEXT = unsafe { nil }
    p_user_data                                voidptr
} 



// VK_EXT_acquire_drm_display is a preprocessor guard. Do not pass it to API calls.
const ext_acquire_drm_display = 1
pub const ext_acquire_drm_display_spec_version = 1
pub const ext_acquire_drm_display_extension_name = "VK_EXT_acquire_drm_display"
type VkAcquireDrmDisplayEXT = fn (     C.PhysicalDevice,     i32,     C.DisplayKHR) Result

pub fn acquire_drm_display_ext(
    physical_device                                 C.PhysicalDevice,
    drm_fd                                          i32,
    display                                         C.DisplayKHR) Result {
      f := VkAcquireDrmDisplayEXT((*loader_p).get_sym('vkAcquireDrmDisplayEXT'
    ) or { 
        println("Couldn't load symbol for 'vkAcquireDrmDisplayEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    drm_fd,
    display)
}


type VkGetDrmDisplayEXT = fn (     C.PhysicalDevice,     i32,     u32,     &C.DisplayKHR) Result

pub fn get_drm_display_ext(
    physical_device                                 C.PhysicalDevice,
    drm_fd                                          i32,
    connector_id                                    u32,
    display                                         &C.DisplayKHR) Result {
      f := VkGetDrmDisplayEXT((*loader_p).get_sym('vkGetDrmDisplayEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetDrmDisplayEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    drm_fd,
    connector_id,
    display)
}




// VK_EXT_robustness2 is a preprocessor guard. Do not pass it to API calls.
const ext_robustness2 = 1
pub const ext_robustness_2_spec_version     = 1
pub const ext_robustness_2_extension_name   = "VK_EXT_robustness2"
// PhysicalDeviceRobustness2FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRobustness2FeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    robust_buffer_access2  Bool32
    robust_image_access2   Bool32
    null_descriptor        Bool32
} 

// PhysicalDeviceRobustness2PropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceRobustness2PropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    robust_storage_buffer_access_size_alignment DeviceSize
    robust_uniform_buffer_access_size_alignment DeviceSize
} 



// VK_EXT_custom_border_color is a preprocessor guard. Do not pass it to API calls.
const ext_custom_border_color = 1
pub const ext_custom_border_color_spec_version = 12
pub const ext_custom_border_color_extension_name = "VK_EXT_custom_border_color"
// SamplerCustomBorderColorCreateInfoEXT extends VkSamplerCreateInfo
pub struct SamplerCustomBorderColorCreateInfoEXT {
mut:
    s_type                   StructureType
    p_next                   voidptr
    custom_border_color      ClearColorValue
    format                   Format
} 

// PhysicalDeviceCustomBorderColorPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceCustomBorderColorPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_custom_border_color_samplers u32
} 

// PhysicalDeviceCustomBorderColorFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceCustomBorderColorFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    custom_border_colors   Bool32
    custom_border_color_without_format Bool32
} 



// VK_GOOGLE_user_type is a preprocessor guard. Do not pass it to API calls.
const google_user_type = 1
pub const google_user_type_spec_version     = 1
pub const google_user_type_extension_name   = "VK_GOOGE_user_type"


// VK_NV_present_barrier is a preprocessor guard. Do not pass it to API calls.
const nv_present_barrier = 1
pub const nv_present_barrier_spec_version   = 1
pub const nv_present_barrier_extension_name = "VK_NV_present_barrier"
// PhysicalDevicePresentBarrierFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePresentBarrierFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    present_barrier        Bool32
} 

// SurfaceCapabilitiesPresentBarrierNV extends VkSurfaceCapabilities2KHR
pub struct SurfaceCapabilitiesPresentBarrierNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    present_barrier_supported Bool32
} 

// SwapchainPresentBarrierCreateInfoNV extends VkSwapchainCreateInfoKHR
pub struct SwapchainPresentBarrierCreateInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    present_barrier_enable Bool32
} 



// VK_EXT_private_data is a preprocessor guard. Do not pass it to API calls.
const ext_private_data = 1
pub const ext_private_data_spec_version     = 1
pub const ext_private_data_extension_name   = "VK_EXT_private_data"
pub type PhysicalDevicePrivateDataFeaturesEXT = PhysicalDevicePrivateDataFeatures

pub type DevicePrivateDataCreateInfoEXT = DevicePrivateDataCreateInfo

pub type PrivateDataSlotCreateInfoEXT = PrivateDataSlotCreateInfo

type VkCreatePrivateDataSlotEXT = fn (     C.Device,     &PrivateDataSlotCreateInfo,     &AllocationCallbacks,     &C.PrivateDataSlot) Result

pub fn create_private_data_slot_ext(
    device                                          C.Device,
    p_create_info                                   &PrivateDataSlotCreateInfo,
    p_allocator                                     &AllocationCallbacks,
    p_private_data_slot                             &C.PrivateDataSlot) Result {
      f := VkCreatePrivateDataSlotEXT((*loader_p).get_sym('vkCreatePrivateDataSlotEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCreatePrivateDataSlotEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_private_data_slot)
}


type VkDestroyPrivateDataSlotEXT = fn (     C.Device,     C.PrivateDataSlot,     &AllocationCallbacks) 

pub fn destroy_private_data_slot_ext(
    device                                          C.Device,
    private_data_slot                               C.PrivateDataSlot,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyPrivateDataSlotEXT((*loader_p).get_sym('vkDestroyPrivateDataSlotEXT'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyPrivateDataSlotEXT': ${err}")
        return 
    })
    f(
    device,
    private_data_slot,
    p_allocator)
}


type VkSetPrivateDataEXT = fn (     C.Device,     ObjectType,     u64,     C.PrivateDataSlot,     u64) Result

pub fn set_private_data_ext(
    device                                          C.Device,
    object_type                                     ObjectType,
    object_handle                                   u64,
    private_data_slot                               C.PrivateDataSlot,
    data                                            u64) Result {
      f := VkSetPrivateDataEXT((*loader_p).get_sym('vkSetPrivateDataEXT'
    ) or { 
        println("Couldn't load symbol for 'vkSetPrivateDataEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    object_type,
    object_handle,
    private_data_slot,
    data)
}


type VkGetPrivateDataEXT = fn (     C.Device,     ObjectType,     u64,     C.PrivateDataSlot,     &u64) 

pub fn get_private_data_ext(
    device                                          C.Device,
    object_type                                     ObjectType,
    object_handle                                   u64,
    private_data_slot                               C.PrivateDataSlot,
    p_data                                          &u64)  {
      f := VkGetPrivateDataEXT((*loader_p).get_sym('vkGetPrivateDataEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetPrivateDataEXT': ${err}")
        return 
    })
    f(
    device,
    object_type,
    object_handle,
    private_data_slot,
    p_data)
}




// VK_EXT_pipeline_creation_cache_control is a preprocessor guard. Do not pass it to API calls.
const ext_pipeline_creation_cache_control = 1
pub const ext_pipeline_creation_cache_control_spec_version = 3
pub const ext_pipeline_creation_cache_control_extension_name = "VK_EXT_pipeline_creation_cache_control"
pub type PhysicalDevicePipelineCreationCacheControlFeaturesEXT = PhysicalDevicePipelineCreationCacheControlFeatures



// VK_NV_device_diagnostics_config is a preprocessor guard. Do not pass it to API calls.
const nv_device_diagnostics_config = 1
pub const nv_device_diagnostics_config_spec_version = 2
pub const nv_device_diagnostics_config_extension_name = "VK_NV_device_diagnostics_config"

pub enum DeviceDiagnosticsConfigFlagBitsNV {
    device_diagnostics_config_enable_shader_debug_info_bit_nv = int(0x00000001)
    device_diagnostics_config_enable_resource_tracking_bit_nv = int(0x00000002)
    device_diagnostics_config_enable_automatic_checkpoints_bit_nv = int(0x00000004)
    device_diagnostics_config_enable_shader_error_reporting_bit_nv = int(0x00000008)
    device_diagnostics_config_flag_bits_max_enum_nv = int(0x7FFFFFFF)
}

pub type DeviceDiagnosticsConfigFlagsNV = u32
// PhysicalDeviceDiagnosticsConfigFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDiagnosticsConfigFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    diagnostics_config     Bool32
} 

// DeviceDiagnosticsConfigCreateInfoNV extends VkDeviceCreateInfo
pub struct DeviceDiagnosticsConfigCreateInfoNV {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    flags                                   DeviceDiagnosticsConfigFlagsNV
} 



// VK_QCOM_render_pass_store_ops is a preprocessor guard. Do not pass it to API calls.
const qcom_render_pass_store_ops = 1
pub const qcom_render_pass_store_ops_spec_version = 2
pub const qcom_render_pass_store_ops_extension_name = "VK_QCOM_render_pass_store_ops"


// VK_NV_cuda_kernel_launch is a preprocessor guard. Do not pass it to API calls.
const nv_cuda_kernel_launch = 1
pub type C.CudaModuleNV = voidptr
pub type C.CudaFunctionNV = voidptr
pub const nv_cuda_kernel_launch_spec_version = 2
pub const nv_cuda_kernel_launch_extension_name = "VK_NV_cuda_kernel_launch"
pub struct CudaModuleCreateInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    data_size              usize
    p_data                 voidptr
} 

pub struct CudaFunctionCreateInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    vkmodule               C.CudaModuleNV
    p_name                 &char
} 

pub struct CudaLaunchInfoNV {
mut:
    s_type                     StructureType
    p_next                     voidptr
    function                   C.CudaFunctionNV
    grid_dim_x                 u32
    grid_dim_y                 u32
    grid_dim_z                 u32
    block_dim_x                u32
    block_dim_y                u32
    block_dim_z                u32
    shared_mem_bytes           u32
    param_count                usize
    p_params                   voidptr
    extra_count                usize
    p_extras                   voidptr
} 

// PhysicalDeviceCudaKernelLaunchFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceCudaKernelLaunchFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    cuda_kernel_launch_features Bool32
} 

// PhysicalDeviceCudaKernelLaunchPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceCudaKernelLaunchPropertiesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    compute_capability_minor u32
    compute_capability_major u32
} 

type VkCreateCudaModuleNV = fn (     C.Device,     &CudaModuleCreateInfoNV,     &AllocationCallbacks,     &C.CudaModuleNV) Result

pub fn create_cuda_module_nv(
    device                                          C.Device,
    p_create_info                                   &CudaModuleCreateInfoNV,
    p_allocator                                     &AllocationCallbacks,
    p_module                                        &C.CudaModuleNV) Result {
      f := VkCreateCudaModuleNV((*loader_p).get_sym('vkCreateCudaModuleNV'
    ) or { 
        println("Couldn't load symbol for 'vkCreateCudaModuleNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_module)
}


type VkGetCudaModuleCacheNV = fn (     C.Device,     C.CudaModuleNV,     &usize,     voidptr) Result

pub fn get_cuda_module_cache_nv(
    device                                          C.Device,
    vkmodule                                        C.CudaModuleNV,
    p_cache_size                                    &usize,
    p_cache_data                                    voidptr) Result {
      f := VkGetCudaModuleCacheNV((*loader_p).get_sym('vkGetCudaModuleCacheNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetCudaModuleCacheNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    vkmodule,
    p_cache_size,
    p_cache_data)
}


type VkCreateCudaFunctionNV = fn (     C.Device,     &CudaFunctionCreateInfoNV,     &AllocationCallbacks,     &C.CudaFunctionNV) Result

pub fn create_cuda_function_nv(
    device                                          C.Device,
    p_create_info                                   &CudaFunctionCreateInfoNV,
    p_allocator                                     &AllocationCallbacks,
    p_function                                      &C.CudaFunctionNV) Result {
      f := VkCreateCudaFunctionNV((*loader_p).get_sym('vkCreateCudaFunctionNV'
    ) or { 
        println("Couldn't load symbol for 'vkCreateCudaFunctionNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_function)
}


type VkDestroyCudaModuleNV = fn (     C.Device,     C.CudaModuleNV,     &AllocationCallbacks) 

pub fn destroy_cuda_module_nv(
    device                                          C.Device,
    vkmodule                                        C.CudaModuleNV,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyCudaModuleNV((*loader_p).get_sym('vkDestroyCudaModuleNV'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyCudaModuleNV': ${err}")
        return 
    })
    f(
    device,
    vkmodule,
    p_allocator)
}


type VkDestroyCudaFunctionNV = fn (     C.Device,     C.CudaFunctionNV,     &AllocationCallbacks) 

pub fn destroy_cuda_function_nv(
    device                                          C.Device,
    function                                        C.CudaFunctionNV,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyCudaFunctionNV((*loader_p).get_sym('vkDestroyCudaFunctionNV'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyCudaFunctionNV': ${err}")
        return 
    })
    f(
    device,
    function,
    p_allocator)
}


type VkCmdCudaLaunchKernelNV = fn (     C.CommandBuffer,     &CudaLaunchInfoNV) 

pub fn cmd_cuda_launch_kernel_nv(
    command_buffer                                  C.CommandBuffer,
    p_launch_info                                   &CudaLaunchInfoNV)  {
      f := VkCmdCudaLaunchKernelNV((*loader_p).get_sym('vkCmdCudaLaunchKernelNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCudaLaunchKernelNV': ${err}")
        return 
    })
    f(
    command_buffer,
    p_launch_info)
}




// VK_NV_low_latency is a preprocessor guard. Do not pass it to API calls.
const nv_low_latency = 1
pub const nv_low_latency_spec_version       = 1
pub const nv_low_latency_extension_name     = "VK_NV_low_latency"
// QueryLowLatencySupportNV extends VkSemaphoreCreateInfo
pub struct QueryLowLatencySupportNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    p_queried_low_latency_data voidptr
} 



// VK_EXT_metal_objects is a preprocessor guard. Do not pass it to API calls.
const ext_metal_objects = 1
pub const ext_metal_objects_spec_version    = 1
pub const ext_metal_objects_extension_name  = "VK_EXT_metal_objects"

pub enum ExportMetalObjectTypeFlagBitsEXT {
    export_metal_object_type_metal_device_bit_ext = int(0x00000001)
    export_metal_object_type_metal_command_queue_bit_ext = int(0x00000002)
    export_metal_object_type_metal_buffer_bit_ext = int(0x00000004)
    export_metal_object_type_metal_texture_bit_ext = int(0x00000008)
    export_metal_object_type_metal_iosurface_bit_ext = int(0x00000010)
    export_metal_object_type_metal_shared_event_bit_ext = int(0x00000020)
    export_metal_object_type_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type ExportMetalObjectTypeFlagsEXT = u32
// ExportMetalObjectCreateInfoEXT extends VkInstanceCreateInfo,VkMemoryAllocateInfo,VkImageCreateInfo,VkImageViewCreateInfo,VkBufferViewCreateInfo,VkSemaphoreCreateInfo,VkEventCreateInfo
pub struct ExportMetalObjectCreateInfoEXT {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    export_object_type                        ExportMetalObjectTypeFlagBitsEXT
} 

pub struct ExportMetalObjectsInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
} 

// ExportMetalDeviceInfoEXT extends VkExportMetalObjectsInfoEXT
pub struct ExportMetalDeviceInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    mtl_device             voidptr
} 

// ExportMetalCommandQueueInfoEXT extends VkExportMetalObjectsInfoEXT
pub struct ExportMetalCommandQueueInfoEXT {
mut:
    s_type                    StructureType
    p_next                    voidptr
    queue                     C.Queue
    mtl_command_queue         voidptr
} 

// ExportMetalBufferInfoEXT extends VkExportMetalObjectsInfoEXT
pub struct ExportMetalBufferInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    memory                 C.DeviceMemory
    mtl_buffer             voidptr
} 

// ImportMetalBufferInfoEXT extends VkMemoryAllocateInfo
pub struct ImportMetalBufferInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    mtl_buffer             voidptr
} 

// ExportMetalTextureInfoEXT extends VkExportMetalObjectsInfoEXT
pub struct ExportMetalTextureInfoEXT {
mut:
    s_type                       StructureType
    p_next                       voidptr
    image                        C.Image
    image_view                   C.ImageView
    buffer_view                  C.BufferView
    plane                        ImageAspectFlagBits
    mtl_texture                  voidptr
} 

// ImportMetalTextureInfoEXT extends VkImageCreateInfo
pub struct ImportMetalTextureInfoEXT {
mut:
    s_type                       StructureType
    p_next                       voidptr
    plane                        ImageAspectFlagBits
    mtl_texture                  voidptr
} 

// ExportMetalIOSurfaceInfoEXT extends VkExportMetalObjectsInfoEXT
pub struct ExportMetalIOSurfaceInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image                  C.Image
    io_surface             voidptr
} 

// ImportMetalIOSurfaceInfoEXT extends VkImageCreateInfo
pub struct ImportMetalIOSurfaceInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    io_surface             voidptr
} 

// ExportMetalSharedEventInfoEXT extends VkExportMetalObjectsInfoEXT
pub struct ExportMetalSharedEventInfoEXT {
mut:
    s_type                   StructureType
    p_next                   voidptr
    semaphore                C.Semaphore
    event                    C.Event
    mtl_shared_event         voidptr
} 

// ImportMetalSharedEventInfoEXT extends VkSemaphoreCreateInfo,VkEventCreateInfo
pub struct ImportMetalSharedEventInfoEXT {
mut:
    s_type                   StructureType
    p_next                   voidptr
    mtl_shared_event         voidptr
} 

type VkExportMetalObjectsEXT = fn (     C.Device,     &ExportMetalObjectsInfoEXT) 

pub fn export_metal_objects_ext(
    device                                          C.Device,
    p_metal_objects_info                            &ExportMetalObjectsInfoEXT)  {
      f := VkExportMetalObjectsEXT((*loader_p).get_sym('vkExportMetalObjectsEXT'
    ) or { 
        println("Couldn't load symbol for 'vkExportMetalObjectsEXT': ${err}")
        return 
    })
    f(
    device,
    p_metal_objects_info)
}




// VK_EXT_descriptor_buffer is a preprocessor guard. Do not pass it to API calls.
const ext_descriptor_buffer = 1
pub type C.AccelerationStructureKHR = voidptr
pub const ext_descriptor_buffer_spec_version = 1
pub const ext_descriptor_buffer_extension_name = "VK_EXT_descriptor_buffer"
// PhysicalDeviceDescriptorBufferPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceDescriptorBufferPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    combined_image_sampler_descriptor_single_array Bool32
    bufferless_push_descriptors Bool32
    allow_sampler_image_view_post_submit_creation Bool32
    descriptor_buffer_offset_alignment DeviceSize
    max_descriptor_buffer_bindings u32
    max_resource_descriptor_buffer_bindings u32
    max_sampler_descriptor_buffer_bindings u32
    max_embedded_immutable_sampler_bindings u32
    max_embedded_immutable_samplers u32
    buffer_capture_replay_descriptor_data_size usize
    image_capture_replay_descriptor_data_size usize
    image_view_capture_replay_descriptor_data_size usize
    sampler_capture_replay_descriptor_data_size usize
    acceleration_structure_capture_replay_descriptor_data_size usize
    sampler_descriptor_size usize
    combined_image_sampler_descriptor_size usize
    sampled_image_descriptor_size usize
    storage_image_descriptor_size usize
    uniform_texel_buffer_descriptor_size usize
    robust_uniform_texel_buffer_descriptor_size usize
    storage_texel_buffer_descriptor_size usize
    robust_storage_texel_buffer_descriptor_size usize
    uniform_buffer_descriptor_size usize
    robust_uniform_buffer_descriptor_size usize
    storage_buffer_descriptor_size usize
    robust_storage_buffer_descriptor_size usize
    input_attachment_descriptor_size usize
    acceleration_structure_descriptor_size usize
    max_sampler_descriptor_buffer_range DeviceSize
    max_resource_descriptor_buffer_range DeviceSize
    sampler_descriptor_buffer_address_space_size DeviceSize
    resource_descriptor_buffer_address_space_size DeviceSize
    descriptor_buffer_address_space_size DeviceSize
} 

// PhysicalDeviceDescriptorBufferDensityMapPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceDescriptorBufferDensityMapPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    combined_image_sampler_density_map_descriptor_size usize
} 

// PhysicalDeviceDescriptorBufferFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDescriptorBufferFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    descriptor_buffer      Bool32
    descriptor_buffer_capture_replay Bool32
    descriptor_buffer_image_layout_ignored Bool32
    descriptor_buffer_push_descriptors Bool32
} 

pub struct DescriptorAddressInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    address                DeviceAddress
    range                  DeviceSize
    format                 Format
} 

pub struct DescriptorBufferBindingInfoEXT {
mut:
    s_type                    StructureType
    p_next                    voidptr
    address                   DeviceAddress
    usage                     BufferUsageFlags
} 

// DescriptorBufferBindingPushDescriptorBufferHandleEXT extends VkDescriptorBufferBindingInfoEXT
pub struct DescriptorBufferBindingPushDescriptorBufferHandleEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    buffer                 C.Buffer
} 

pub union DescriptorDataEXT {
mut:
    p_sampler                                &C.Sampler
    p_combined_image_sampler                 &DescriptorImageInfo
    p_input_attachment_image                 &DescriptorImageInfo
    p_sampled_image                          &DescriptorImageInfo
    p_storage_image                          &DescriptorImageInfo
    p_uniform_texel_buffer                   &DescriptorAddressInfoEXT
    p_storage_texel_buffer                   &DescriptorAddressInfoEXT
    p_uniform_buffer                         &DescriptorAddressInfoEXT
    p_storage_buffer                         &DescriptorAddressInfoEXT
    acceleration_structure                   DeviceAddress
} 

pub struct DescriptorGetInfoEXT {
mut:
    s_type                     StructureType
    p_next                     voidptr
    vktype                     DescriptorType
    data                       DescriptorDataEXT
} 

pub struct BufferCaptureDescriptorDataInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    buffer                 C.Buffer
} 

pub struct ImageCaptureDescriptorDataInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image                  C.Image
} 

pub struct ImageViewCaptureDescriptorDataInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image_view             C.ImageView
} 

pub struct SamplerCaptureDescriptorDataInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    sampler                C.Sampler
} 

// OpaqueCaptureDescriptorDataCreateInfoEXT extends VkBufferCreateInfo,VkImageCreateInfo,VkImageViewCreateInfo,VkSamplerCreateInfo,VkAccelerationStructureCreateInfoKHR,VkAccelerationStructureCreateInfoNV
pub struct OpaqueCaptureDescriptorDataCreateInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    opaque_capture_descriptor_data voidptr
} 

pub struct AccelerationStructureCaptureDescriptorDataInfoEXT {
mut:
    s_type                            StructureType
    p_next                            voidptr
    acceleration_structure            C.AccelerationStructureKHR
    acceleration_structure_nv         C.AccelerationStructureNV
} 

type VkGetDescriptorSetLayoutSizeEXT = fn (     C.Device,     C.DescriptorSetLayout,     &DeviceSize) 

pub fn get_descriptor_set_layout_size_ext(
    device                                          C.Device,
    layout                                          C.DescriptorSetLayout,
    p_layout_size_in_bytes                          &DeviceSize)  {
      f := VkGetDescriptorSetLayoutSizeEXT((*loader_p).get_sym('vkGetDescriptorSetLayoutSizeEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetDescriptorSetLayoutSizeEXT': ${err}")
        return 
    })
    f(
    device,
    layout,
    p_layout_size_in_bytes)
}


type VkGetDescriptorSetLayoutBindingOffsetEXT = fn (     C.Device,     C.DescriptorSetLayout,     u32,     &DeviceSize) 

pub fn get_descriptor_set_layout_binding_offset_ext(
    device                                          C.Device,
    layout                                          C.DescriptorSetLayout,
    binding                                         u32,
    p_offset                                        &DeviceSize)  {
      f := VkGetDescriptorSetLayoutBindingOffsetEXT((*loader_p).get_sym('vkGetDescriptorSetLayoutBindingOffsetEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetDescriptorSetLayoutBindingOffsetEXT': ${err}")
        return 
    })
    f(
    device,
    layout,
    binding,
    p_offset)
}


type VkGetDescriptorEXT = fn (     C.Device,     &DescriptorGetInfoEXT,     usize,     voidptr) 

pub fn get_descriptor_ext(
    device                                          C.Device,
    p_descriptor_info                               &DescriptorGetInfoEXT,
    data_size                                       usize,
    p_descriptor                                    voidptr)  {
      f := VkGetDescriptorEXT((*loader_p).get_sym('vkGetDescriptorEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetDescriptorEXT': ${err}")
        return 
    })
    f(
    device,
    p_descriptor_info,
    data_size,
    p_descriptor)
}


type VkCmdBindDescriptorBuffersEXT = fn (     C.CommandBuffer,     u32,     &DescriptorBufferBindingInfoEXT) 

pub fn cmd_bind_descriptor_buffers_ext(
    command_buffer                                  C.CommandBuffer,
    buffer_count                                    u32,
    p_binding_infos                                 &DescriptorBufferBindingInfoEXT)  {
      f := VkCmdBindDescriptorBuffersEXT((*loader_p).get_sym('vkCmdBindDescriptorBuffersEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindDescriptorBuffersEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer_count,
    p_binding_infos)
}


type VkCmdSetDescriptorBufferOffsetsEXT = fn (     C.CommandBuffer,     PipelineBindPoint,     C.PipelineLayout,     u32,     u32,     &u32,     &DeviceSize) 

pub fn cmd_set_descriptor_buffer_offsets_ext(
    command_buffer                                  C.CommandBuffer,
    pipeline_bind_point                             PipelineBindPoint,
    layout                                          C.PipelineLayout,
    first_set                                       u32,
    set_count                                       u32,
    p_buffer_indices                                &u32,
    p_offsets                                       &DeviceSize)  {
      f := VkCmdSetDescriptorBufferOffsetsEXT((*loader_p).get_sym('vkCmdSetDescriptorBufferOffsetsEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDescriptorBufferOffsetsEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    pipeline_bind_point,
    layout,
    first_set,
    set_count,
    p_buffer_indices,
    p_offsets)
}


type VkCmdBindDescriptorBufferEmbeddedSamplersEXT = fn (     C.CommandBuffer,     PipelineBindPoint,     C.PipelineLayout,     u32) 

pub fn cmd_bind_descriptor_buffer_embedded_samplers_ext(
    command_buffer                                  C.CommandBuffer,
    pipeline_bind_point                             PipelineBindPoint,
    layout                                          C.PipelineLayout,
    set                                             u32)  {
      f := VkCmdBindDescriptorBufferEmbeddedSamplersEXT((*loader_p).get_sym('vkCmdBindDescriptorBufferEmbeddedSamplersEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindDescriptorBufferEmbeddedSamplersEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    pipeline_bind_point,
    layout,
    set)
}


type VkGetBufferOpaqueCaptureDescriptorDataEXT = fn (     C.Device,     &BufferCaptureDescriptorDataInfoEXT,     voidptr) Result

pub fn get_buffer_opaque_capture_descriptor_data_ext(
    device                                          C.Device,
    p_info                                          &BufferCaptureDescriptorDataInfoEXT,
    p_data                                          voidptr) Result {
      f := VkGetBufferOpaqueCaptureDescriptorDataEXT((*loader_p).get_sym('vkGetBufferOpaqueCaptureDescriptorDataEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetBufferOpaqueCaptureDescriptorDataEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_info,
    p_data)
}


type VkGetImageOpaqueCaptureDescriptorDataEXT = fn (     C.Device,     &ImageCaptureDescriptorDataInfoEXT,     voidptr) Result

pub fn get_image_opaque_capture_descriptor_data_ext(
    device                                          C.Device,
    p_info                                          &ImageCaptureDescriptorDataInfoEXT,
    p_data                                          voidptr) Result {
      f := VkGetImageOpaqueCaptureDescriptorDataEXT((*loader_p).get_sym('vkGetImageOpaqueCaptureDescriptorDataEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageOpaqueCaptureDescriptorDataEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_info,
    p_data)
}


type VkGetImageViewOpaqueCaptureDescriptorDataEXT = fn (     C.Device,     &ImageViewCaptureDescriptorDataInfoEXT,     voidptr) Result

pub fn get_image_view_opaque_capture_descriptor_data_ext(
    device                                          C.Device,
    p_info                                          &ImageViewCaptureDescriptorDataInfoEXT,
    p_data                                          voidptr) Result {
      f := VkGetImageViewOpaqueCaptureDescriptorDataEXT((*loader_p).get_sym('vkGetImageViewOpaqueCaptureDescriptorDataEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetImageViewOpaqueCaptureDescriptorDataEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_info,
    p_data)
}


type VkGetSamplerOpaqueCaptureDescriptorDataEXT = fn (     C.Device,     &SamplerCaptureDescriptorDataInfoEXT,     voidptr) Result

pub fn get_sampler_opaque_capture_descriptor_data_ext(
    device                                          C.Device,
    p_info                                          &SamplerCaptureDescriptorDataInfoEXT,
    p_data                                          voidptr) Result {
      f := VkGetSamplerOpaqueCaptureDescriptorDataEXT((*loader_p).get_sym('vkGetSamplerOpaqueCaptureDescriptorDataEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetSamplerOpaqueCaptureDescriptorDataEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_info,
    p_data)
}


type VkGetAccelerationStructureOpaqueCaptureDescriptorDataEXT = fn (     C.Device,     &AccelerationStructureCaptureDescriptorDataInfoEXT,     voidptr) Result

pub fn get_acceleration_structure_opaque_capture_descriptor_data_ext(
    device                                          C.Device,
    p_info                                          &AccelerationStructureCaptureDescriptorDataInfoEXT,
    p_data                                          voidptr) Result {
      f := VkGetAccelerationStructureOpaqueCaptureDescriptorDataEXT((*loader_p).get_sym('vkGetAccelerationStructureOpaqueCaptureDescriptorDataEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetAccelerationStructureOpaqueCaptureDescriptorDataEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_info,
    p_data)
}




// VK_EXT_graphics_pipeline_library is a preprocessor guard. Do not pass it to API calls.
const ext_graphics_pipeline_library = 1
pub const ext_graphics_pipeline_library_spec_version = 1
pub const ext_graphics_pipeline_library_extension_name = "VK_EXT_graphics_pipeline_library"

pub enum GraphicsPipelineLibraryFlagBitsEXT {
    graphics_pipeline_library_vertex_input_interface_bit_ext = int(0x00000001)
    graphics_pipeline_library_pre_rasterization_shaders_bit_ext = int(0x00000002)
    graphics_pipeline_library_fragment_shader_bit_ext = int(0x00000004)
    graphics_pipeline_library_fragment_output_interface_bit_ext = int(0x00000008)
    graphics_pipeline_library_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type GraphicsPipelineLibraryFlagsEXT = u32
// PhysicalDeviceGraphicsPipelineLibraryFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceGraphicsPipelineLibraryFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    graphics_pipeline_library Bool32
} 

// PhysicalDeviceGraphicsPipelineLibraryPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceGraphicsPipelineLibraryPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    graphics_pipeline_library_fast_linking Bool32
    graphics_pipeline_library_independent_interpolation_decoration Bool32
} 

// GraphicsPipelineLibraryCreateInfoEXT extends VkGraphicsPipelineCreateInfo
pub struct GraphicsPipelineLibraryCreateInfoEXT {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    flags                                    GraphicsPipelineLibraryFlagsEXT
} 



// VK_AMD_shader_early_and_late_fragment_tests is a preprocessor guard. Do not pass it to API calls.
const amd_shader_early_and_late_fragment_tests = 1
pub const amd_shader_early_and_late_fragment_tests_spec_version = 1
pub const amd_shader_early_and_late_fragment_tests_extension_name = "VK_AMD_shader_early_and_late_fragment_tests"
// PhysicalDeviceShaderEarlyAndLateFragmentTestsFeaturesAMD extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderEarlyAndLateFragmentTestsFeaturesAMD {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_early_and_late_fragment_tests Bool32
} 



// VK_NV_fragment_shading_rate_enums is a preprocessor guard. Do not pass it to API calls.
const nv_fragment_shading_rate_enums = 1
pub const nv_fragment_shading_rate_enums_spec_version = 1
pub const nv_fragment_shading_rate_enums_extension_name = "VK_NV_fragment_shading_rate_enums"

pub enum FragmentShadingRateTypeNV {
    fragment_shading_rate_type_fragment_size_nv = int(0)
    fragment_shading_rate_type_enums_nv = int(1)
    fragment_shading_rate_type_max_enum_nv = int(0x7FFFFFFF)
}


pub enum FragmentShadingRateNV {
    fragment_shading_rate_1_invocation_per_pixel_nv = int(0)
    fragment_shading_rate_1_invocation_per_1x2_pixels_nv = int(1)
    fragment_shading_rate_1_invocation_per_2x1_pixels_nv = int(4)
    fragment_shading_rate_1_invocation_per_2x2_pixels_nv = int(5)
    fragment_shading_rate_1_invocation_per_2x4_pixels_nv = int(6)
    fragment_shading_rate_1_invocation_per_4x2_pixels_nv = int(9)
    fragment_shading_rate_1_invocation_per_4x4_pixels_nv = int(10)
    fragment_shading_rate_2_invocations_per_pixel_nv = int(11)
    fragment_shading_rate_4_invocations_per_pixel_nv = int(12)
    fragment_shading_rate_8_invocations_per_pixel_nv = int(13)
    fragment_shading_rate_16_invocations_per_pixel_nv = int(14)
    fragment_shading_rate_no_invocations_nv = int(15)
    fragment_shading_rate_max_enum_nv = int(0x7FFFFFFF)
}

// PhysicalDeviceFragmentShadingRateEnumsFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceFragmentShadingRateEnumsFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    fragment_shading_rate_enums Bool32
    supersample_fragment_shading_rates Bool32
    no_invocation_fragment_shading_rates Bool32
} 

// PhysicalDeviceFragmentShadingRateEnumsPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceFragmentShadingRateEnumsPropertiesNV {
mut:
    s_type                       StructureType
    p_next                       voidptr
    max_fragment_shading_rate_invocation_count SampleCountFlagBits
} 

// PipelineFragmentShadingRateEnumStateCreateInfoNV extends VkGraphicsPipelineCreateInfo
pub struct PipelineFragmentShadingRateEnumStateCreateInfoNV {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    shading_rate_type                         FragmentShadingRateTypeNV
    shading_rate                              FragmentShadingRateNV
    combiner_ops                              []FragmentShadingRateCombinerOpKHR
} 

type VkCmdSetFragmentShadingRateEnumNV = fn (     C.CommandBuffer,     FragmentShadingRateNV,     []FragmentShadingRateCombinerOpKHR) 

pub fn cmd_set_fragment_shading_rate_enum_nv(
    command_buffer                                  C.CommandBuffer,
    shading_rate                                    FragmentShadingRateNV,
    combiner_ops                                    []FragmentShadingRateCombinerOpKHR)  {
      f := VkCmdSetFragmentShadingRateEnumNV((*loader_p).get_sym('vkCmdSetFragmentShadingRateEnumNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetFragmentShadingRateEnumNV': ${err}")
        return 
    })
    f(
    command_buffer,
    shading_rate,
    combiner_ops)
}




// VK_NV_ray_tracing_motion_blur is a preprocessor guard. Do not pass it to API calls.
const nv_ray_tracing_motion_blur = 1
pub const nv_ray_tracing_motion_blur_spec_version = 1
pub const nv_ray_tracing_motion_blur_extension_name = "VK_NV_ray_tracing_motion_blur"

pub enum AccelerationStructureMotionInstanceTypeNV {
    acceleration_structure_motion_instance_type_static_nv = int(0)
    acceleration_structure_motion_instance_type_matrix_motion_nv = int(1)
    acceleration_structure_motion_instance_type_srt_motion_nv = int(2)
    acceleration_structure_motion_instance_type_max_enum_nv = int(0x7FFFFFFF)
}

pub type AccelerationStructureMotionInfoFlagsNV = u32
pub type AccelerationStructureMotionInstanceFlagsNV = u32
pub union DeviceOrHostAddressConstKHR {
mut:
    device_address         DeviceAddress
    host_address           voidptr
} 

// AccelerationStructureGeometryMotionTrianglesDataNV extends VkAccelerationStructureGeometryTrianglesDataKHR
pub struct AccelerationStructureGeometryMotionTrianglesDataNV {
mut:
    s_type                               StructureType
    p_next                               voidptr
    vertex_data                          DeviceOrHostAddressConstKHR
} 

// AccelerationStructureMotionInfoNV extends VkAccelerationStructureCreateInfoKHR
pub struct AccelerationStructureMotionInfoNV {
mut:
    s_type                                          StructureType
    p_next                                          voidptr
    max_instances                                   u32
    flags                                           AccelerationStructureMotionInfoFlagsNV
} 

pub struct AccelerationStructureMatrixMotionInstanceNV {
mut:
    transform_t0                      TransformMatrixKHR
    transform_t1                      TransformMatrixKHR
    instance_custom_index             u32
    mask                              u32
    instance_shader_binding_table_record_offset u32
    flags                             GeometryInstanceFlagsKHR
    acceleration_structure_reference  u64
} 

pub struct SRTDataNV {
mut:
    sx           f32
    a            f32
    b            f32
    pvx          f32
    sy           f32
    c            f32
    pvy          f32
    sz           f32
    pvz          f32
    qx           f32
    qy           f32
    qz           f32
    qw           f32
    tx           f32
    ty           f32
    tz           f32
} 

pub struct AccelerationStructureSRTMotionInstanceNV {
mut:
    transform_t0                      SRTDataNV
    transform_t1                      SRTDataNV
    instance_custom_index             u32
    mask                              u32
    instance_shader_binding_table_record_offset u32
    flags                             GeometryInstanceFlagsKHR
    acceleration_structure_reference  u64
} 

pub union AccelerationStructureMotionInstanceDataNV {
mut:
    static_instance                                      AccelerationStructureInstanceKHR
    matrix_motion_instance                               AccelerationStructureMatrixMotionInstanceNV
    srt_motion_instance                                  AccelerationStructureSRTMotionInstanceNV
} 

pub struct AccelerationStructureMotionInstanceNV {
mut:
    vktype                                              AccelerationStructureMotionInstanceTypeNV
    flags                                               AccelerationStructureMotionInstanceFlagsNV
    data                                                AccelerationStructureMotionInstanceDataNV
} 

// PhysicalDeviceRayTracingMotionBlurFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRayTracingMotionBlurFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    ray_tracing_motion_blur Bool32
    ray_tracing_motion_blur_pipeline_trace_rays_indirect Bool32
} 



// VK_EXT_ycbcr_2plane_444_formats is a preprocessor guard. Do not pass it to API calls.
const ext_ycbcr_2plane_444_formats = 1
pub const ext_ycbcr_2plane_444_formats_spec_version = 1
pub const ext_ycbcr_2plane_444_formats_extension_name = "VK_EXT_ycbcr_2plane_444_formats"
// PhysicalDeviceYcbcr2Plane444FormatsFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceYcbcr2Plane444FormatsFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    ycbcr2plane444_formats Bool32
} 



// VK_EXT_fragment_density_map2 is a preprocessor guard. Do not pass it to API calls.
const ext_fragment_density_map2 = 1
pub const ext_fragment_density_map_2_spec_version = 1
pub const ext_fragment_density_map_2_extension_name = "VK_EXT_fragment_density_map2"
// PhysicalDeviceFragmentDensityMap2FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceFragmentDensityMap2FeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    fragment_density_map_deferred Bool32
} 

// PhysicalDeviceFragmentDensityMap2PropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceFragmentDensityMap2PropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    subsampled_loads       Bool32
    subsampled_coarse_reconstruction_early_access Bool32
    max_subsampled_array_layers u32
    max_descriptor_set_subsampled_samplers u32
} 



// VK_QCOM_rotated_copy_commands is a preprocessor guard. Do not pass it to API calls.
const qcom_rotated_copy_commands = 1
pub const qcom_rotated_copy_commands_spec_version = 1
pub const qcom_rotated_copy_commands_extension_name = "VK_QCOM_rotated_copy_commands"
// CopyCommandTransformInfoQCOM extends VkBufferImageCopy2,VkImageBlit2
pub struct CopyCommandTransformInfoQCOM {
mut:
    s_type                               StructureType
    p_next                               voidptr
    transform                            SurfaceTransformFlagBitsKHR
} 



// VK_EXT_image_robustness is a preprocessor guard. Do not pass it to API calls.
const ext_image_robustness = 1
pub const ext_image_robustness_spec_version = 1
pub const ext_image_robustness_extension_name = "VK_EXT_image_robustness"
pub type PhysicalDeviceImageRobustnessFeaturesEXT = PhysicalDeviceImageRobustnessFeatures



// VK_EXT_image_compression_control is a preprocessor guard. Do not pass it to API calls.
const ext_image_compression_control = 1
pub const ext_image_compression_control_spec_version = 1
pub const ext_image_compression_control_extension_name = "VK_EXT_image_compression_control"

pub enum ImageCompressionFlagBitsEXT {
    image_compression_default_ext = int(0)
    image_compression_fixed_rate_default_ext = int(0x00000001)
    image_compression_fixed_rate_explicit_ext = int(0x00000002)
    image_compression_disabled_ext = int(0x00000004)
    image_compression_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type ImageCompressionFlagsEXT = u32

pub enum ImageCompressionFixedRateFlagBitsEXT {
    image_compression_fixed_rate_none_ext = int(0)
    image_compression_fixed_rate_1bpc_bit_ext = int(0x00000001)
    image_compression_fixed_rate_2bpc_bit_ext = int(0x00000002)
    image_compression_fixed_rate_3bpc_bit_ext = int(0x00000004)
    image_compression_fixed_rate_4bpc_bit_ext = int(0x00000008)
    image_compression_fixed_rate_5bpc_bit_ext = int(0x00000010)
    image_compression_fixed_rate_6bpc_bit_ext = int(0x00000020)
    image_compression_fixed_rate_7bpc_bit_ext = int(0x00000040)
    image_compression_fixed_rate_8bpc_bit_ext = int(0x00000080)
    image_compression_fixed_rate_9bpc_bit_ext = int(0x00000100)
    image_compression_fixed_rate_10bpc_bit_ext = int(0x00000200)
    image_compression_fixed_rate_11bpc_bit_ext = int(0x00000400)
    image_compression_fixed_rate_12bpc_bit_ext = int(0x00000800)
    image_compression_fixed_rate_13bpc_bit_ext = int(0x00001000)
    image_compression_fixed_rate_14bpc_bit_ext = int(0x00002000)
    image_compression_fixed_rate_15bpc_bit_ext = int(0x00004000)
    image_compression_fixed_rate_16bpc_bit_ext = int(0x00008000)
    image_compression_fixed_rate_17bpc_bit_ext = int(0x00010000)
    image_compression_fixed_rate_18bpc_bit_ext = int(0x00020000)
    image_compression_fixed_rate_19bpc_bit_ext = int(0x00040000)
    image_compression_fixed_rate_20bpc_bit_ext = int(0x00080000)
    image_compression_fixed_rate_21bpc_bit_ext = int(0x00100000)
    image_compression_fixed_rate_22bpc_bit_ext = int(0x00200000)
    image_compression_fixed_rate_23bpc_bit_ext = int(0x00400000)
    image_compression_fixed_rate_24bpc_bit_ext = int(0x00800000)
    image_compression_fixed_rate_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type ImageCompressionFixedRateFlagsEXT = u32
// PhysicalDeviceImageCompressionControlFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceImageCompressionControlFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image_compression_control Bool32
} 

// ImageCompressionControlEXT extends VkImageCreateInfo,VkSwapchainCreateInfoKHR,VkPhysicalDeviceImageFormatInfo2
pub struct ImageCompressionControlEXT {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    flags                                       ImageCompressionFlagsEXT
    compression_control_plane_count             u32
    p_fixed_rate_flags                          &ImageCompressionFixedRateFlagsEXT
} 

// ImageCompressionPropertiesEXT extends VkImageFormatProperties2,VkSurfaceFormat2KHR,VkSubresourceLayout2KHR
pub struct ImageCompressionPropertiesEXT {
mut:
    s_type                                     StructureType
    p_next                                     voidptr
    image_compression_flags                    ImageCompressionFlagsEXT
    image_compression_fixed_rate_flags         ImageCompressionFixedRateFlagsEXT
} 



// VK_EXT_attachment_feedback_loop_layout is a preprocessor guard. Do not pass it to API calls.
const ext_attachment_feedback_loop_layout = 1
pub const ext_attachment_feedback_loop_layout_spec_version = 2
pub const ext_attachment_feedback_loop_layout_extension_name = "VK_EXT_attachment_feedback_loop_layout"
// PhysicalDeviceAttachmentFeedbackLoopLayoutFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceAttachmentFeedbackLoopLayoutFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    attachment_feedback_loop_layout Bool32
} 



// VK_EXT_4444_formats is a preprocessor guard. Do not pass it to API calls.
const ext_4444_formats = 1
pub const ext_4444_formats_spec_version     = 1
pub const ext_4444_formats_extension_name   = "VK_EXT_4444_formats"
// PhysicalDevice4444FormatsFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevice4444FormatsFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    format_a4_r4_g4_b4     Bool32
    format_a4_b4_g4_r4     Bool32
} 



// VK_EXT_device_fault is a preprocessor guard. Do not pass it to API calls.
const ext_device_fault = 1
pub const ext_device_fault_spec_version     = 2
pub const ext_device_fault_extension_name   = "VK_EXT_device_fault"

pub enum DeviceFaultAddressTypeEXT {
    device_fault_address_type_none_ext = int(0)
    device_fault_address_type_read_invalid_ext = int(1)
    device_fault_address_type_write_invalid_ext = int(2)
    device_fault_address_type_execute_invalid_ext = int(3)
    device_fault_address_type_instruction_pointer_unknown_ext = int(4)
    device_fault_address_type_instruction_pointer_invalid_ext = int(5)
    device_fault_address_type_instruction_pointer_fault_ext = int(6)
    device_fault_address_type_max_enum_ext = int(0x7FFFFFFF)
}


pub enum DeviceFaultVendorBinaryHeaderVersionEXT {
    device_fault_vendor_binary_header_version_one_ext = int(1)
    device_fault_vendor_binary_header_version_max_enum_ext = int(0x7FFFFFFF)
}

// PhysicalDeviceFaultFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceFaultFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_fault           Bool32
    device_fault_vendor_binary Bool32
} 

pub struct DeviceFaultCountsEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    address_info_count     u32
    vendor_info_count      u32
    vendor_binary_size     DeviceSize
} 

pub struct DeviceFaultAddressInfoEXT {
mut:
    address_type                       DeviceFaultAddressTypeEXT
    reported_address                   DeviceAddress
    address_precision                  DeviceSize
} 

pub struct DeviceFaultVendorInfoEXT {
mut:
    description     []char
    vendor_fault_code u64
    vendor_fault_data u64
} 

pub struct DeviceFaultInfoEXT {
mut:
    s_type                              StructureType
    p_next                              voidptr
    description                         []char
    p_address_infos                     &DeviceFaultAddressInfoEXT
    p_vendor_infos                      &DeviceFaultVendorInfoEXT
    p_vendor_binary_data                voidptr
} 

pub struct DeviceFaultVendorBinaryHeaderVersionOneEXT {
mut:
    header_size                                      u32
    header_version                                   DeviceFaultVendorBinaryHeaderVersionEXT
    vendor_id                                        u32
    device_id                                        u32
    driver_version                                   u32
    pipeline_cache_uuid                              []u8
    application_name_offset                          u32
    application_version                              u32
    engine_name_offset                               u32
    engine_version                                   u32
    api_version                                      u32
} 

type VkGetDeviceFaultInfoEXT = fn (     C.Device,     &DeviceFaultCountsEXT,     &DeviceFaultInfoEXT) Result

pub fn get_device_fault_info_ext(
    device                                          C.Device,
    p_fault_counts                                  &DeviceFaultCountsEXT,
    p_fault_info                                    &DeviceFaultInfoEXT) Result {
      f := VkGetDeviceFaultInfoEXT((*loader_p).get_sym('vkGetDeviceFaultInfoEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceFaultInfoEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_fault_counts,
    p_fault_info)
}




// VK_ARM_rasterization_order_attachment_access is a preprocessor guard. Do not pass it to API calls.
const arm_rasterization_order_attachment_access = 1
pub const arm_rasterization_order_attachment_access_spec_version = 1
pub const arm_rasterization_order_attachment_access_extension_name = "VK_ARM_rasterization_order_attachment_access"
// PhysicalDeviceRasterizationOrderAttachmentAccessFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRasterizationOrderAttachmentAccessFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    rasterization_order_color_attachment_access Bool32
    rasterization_order_depth_attachment_access Bool32
    rasterization_order_stencil_attachment_access Bool32
} 

pub type PhysicalDeviceRasterizationOrderAttachmentAccessFeaturesARM = PhysicalDeviceRasterizationOrderAttachmentAccessFeaturesEXT



// VK_EXT_rgba10x6_formats is a preprocessor guard. Do not pass it to API calls.
const ext_rgba10x6_formats = 1
pub const ext_rgba10x6_formats_spec_version = 1
pub const ext_rgba10x6_formats_extension_name = "VK_EXT_rgba10x6_formats"
// PhysicalDeviceRGBA10X6FormatsFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRGBA10X6FormatsFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    format_rgba10x6_without_y_cb_cr_sampler Bool32
} 



// VK_NV_acquire_winrt_display is a preprocessor guard. Do not pass it to API calls.
const nv_acquire_winrt_display = 1
pub const nv_acquire_winrt_display_spec_version = 1
pub const nv_acquire_winrt_display_extension_name = "VK_NV_acquire_winrt_display"
type VkAcquireWinrtDisplayNV = fn (     C.PhysicalDevice,     C.DisplayKHR) Result

pub fn acquire_winrt_display_nv(
    physical_device                                 C.PhysicalDevice,
    display                                         C.DisplayKHR) Result {
      f := VkAcquireWinrtDisplayNV((*loader_p).get_sym('vkAcquireWinrtDisplayNV'
    ) or { 
        println("Couldn't load symbol for 'vkAcquireWinrtDisplayNV': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    display)
}


type VkGetWinrtDisplayNV = fn (     C.PhysicalDevice,     u32,     &C.DisplayKHR) Result

pub fn get_winrt_display_nv(
    physical_device                                 C.PhysicalDevice,
    device_relative_id                              u32,
    p_display                                       &C.DisplayKHR) Result {
      f := VkGetWinrtDisplayNV((*loader_p).get_sym('vkGetWinrtDisplayNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetWinrtDisplayNV': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    device_relative_id,
    p_display)
}




// VK_EXT_directfb_surface is a preprocessor guard. Do not pass it to API calls.
const ext_directfb_surface = 1
pub const ext_directfb_surface_spec_version = 1
pub const ext_directfb_surface_extension_name = "VK_EXT_directfb_surface"
pub type DirectFBSurfaceCreateFlagsEXT = u32
pub struct DirectFBSurfaceCreateInfoEXT {
mut:
    s_type                                 StructureType
    p_next                                 voidptr
    flags                                  DirectFBSurfaceCreateFlagsEXT
    dfb                                    voidptr
    surface                                voidptr
} 

type VkCreateDirectFBSurfaceEXT = fn (     C.Instance,     &DirectFBSurfaceCreateInfoEXT,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_direct_fb_surface_ext(
    instance                                        C.Instance,
    p_create_info                                   &DirectFBSurfaceCreateInfoEXT,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateDirectFBSurfaceEXT((*loader_p).get_sym('vkCreateDirectFBSurfaceEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCreateDirectFBSurfaceEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}


type VkGetPhysicalDeviceDirectFBPresentationSupportEXT = fn (     C.PhysicalDevice,     u32,     voidptr) Bool32

pub fn get_physical_device_direct_fb_presentation_support_ext(
    physical_device                                 C.PhysicalDevice,
    queue_family_index                              u32,
    dfb                                             voidptr) Bool32 {
      f := VkGetPhysicalDeviceDirectFBPresentationSupportEXT((*loader_p).get_sym("vkGetPhysicalDeviceDirectFBPresentationSupportEXT"
    ) or { 
        panic("Couldn't load symbol for 'vkGetPhysicalDeviceDirectFBPresentationSupportEXT': ${err}") })
    return f(
    physical_device,
    queue_family_index,
    dfb)
}




// VK_VALVE_mutable_descriptor_type is a preprocessor guard. Do not pass it to API calls.
const valve_mutable_descriptor_type = 1
pub const valve_mutable_descriptor_type_spec_version = 1
pub const valve_mutable_descriptor_type_extension_name = "VK_VAVE_mutable_descriptor_type"
// PhysicalDeviceMutableDescriptorTypeFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMutableDescriptorTypeFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    mutable_descriptor_type Bool32
} 

pub type PhysicalDeviceMutableDescriptorTypeFeaturesVALVE = PhysicalDeviceMutableDescriptorTypeFeaturesEXT

pub struct MutableDescriptorTypeListEXT {
mut:
    descriptor_type_count          u32
    p_descriptor_types             &DescriptorType
} 

pub type MutableDescriptorTypeListVALVE = MutableDescriptorTypeListEXT

// MutableDescriptorTypeCreateInfoEXT extends VkDescriptorSetLayoutCreateInfo,VkDescriptorPoolCreateInfo
pub struct MutableDescriptorTypeCreateInfoEXT {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    mutable_descriptor_type_list_count           u32
    p_mutable_descriptor_type_lists              &MutableDescriptorTypeListEXT
} 

pub type MutableDescriptorTypeCreateInfoVALVE = MutableDescriptorTypeCreateInfoEXT



// VK_EXT_vertex_input_dynamic_state is a preprocessor guard. Do not pass it to API calls.
const ext_vertex_input_dynamic_state = 1
pub const ext_vertex_input_dynamic_state_spec_version = 2
pub const ext_vertex_input_dynamic_state_extension_name = "VK_EXT_vertex_input_dynamic_state"
// PhysicalDeviceVertexInputDynamicStateFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceVertexInputDynamicStateFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    vertex_input_dynamic_state Bool32
} 

pub struct VertexInputBindingDescription2EXT {
mut:
    s_type                   StructureType
    p_next                   voidptr
    binding                  u32
    stride                   u32
    input_rate               VertexInputRate
    divisor                  u32
} 

pub struct VertexInputAttributeDescription2EXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    location               u32
    binding                u32
    format                 Format
    offset                 u32
} 

type VkCmdSetVertexInputEXT = fn (     C.CommandBuffer,     u32,     &VertexInputBindingDescription2EXT,     u32,     &VertexInputAttributeDescription2EXT) 

pub fn cmd_set_vertex_input_ext(
    command_buffer                                  C.CommandBuffer,
    vertex_binding_description_count                u32,
    p_vertex_binding_descriptions                   &VertexInputBindingDescription2EXT,
    vertex_attribute_description_count              u32,
    p_vertex_attribute_descriptions                 &VertexInputAttributeDescription2EXT)  {
      f := VkCmdSetVertexInputEXT((*loader_p).get_sym('vkCmdSetVertexInputEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetVertexInputEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    vertex_binding_description_count,
    p_vertex_binding_descriptions,
    vertex_attribute_description_count,
    p_vertex_attribute_descriptions)
}




// VK_EXT_physical_device_drm is a preprocessor guard. Do not pass it to API calls.
const ext_physical_device_drm = 1
pub const ext_physical_device_drm_spec_version = 1
pub const ext_physical_device_drm_extension_name = "VK_EXT_physical_device_drm"
// PhysicalDeviceDrmPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceDrmPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    has_primary            Bool32
    has_render             Bool32
    primary_major          i64
    primary_minor          i64
    render_major           i64
    render_minor           i64
} 



// VK_EXT_device_address_binding_report is a preprocessor guard. Do not pass it to API calls.
const ext_device_address_binding_report = 1
pub const ext_device_address_binding_report_spec_version = 1
pub const ext_device_address_binding_report_extension_name = "VK_EXT_device_address_binding_report"

pub enum DeviceAddressBindingTypeEXT {
    device_address_binding_type_bind_ext = int(0)
    device_address_binding_type_unbind_ext = int(1)
    device_address_binding_type_max_enum_ext = int(0x7FFFFFFF)
}


pub enum DeviceAddressBindingFlagBitsEXT {
    device_address_binding_internal_object_bit_ext = int(0x00000001)
    device_address_binding_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type DeviceAddressBindingFlagsEXT = u32
// PhysicalDeviceAddressBindingReportFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceAddressBindingReportFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    report_address_binding Bool32
} 

// DeviceAddressBindingCallbackDataEXT extends VkDebugUtilsMessengerCallbackDataEXT
pub struct DeviceAddressBindingCallbackDataEXT {
mut:
    s_type                                StructureType
    p_next                                voidptr
    flags                                 DeviceAddressBindingFlagsEXT
    base_address                          DeviceAddress
    size                                  DeviceSize
    binding_type                          DeviceAddressBindingTypeEXT
} 



// VK_EXT_depth_clip_control is a preprocessor guard. Do not pass it to API calls.
const ext_depth_clip_control = 1
pub const ext_depth_clip_control_spec_version = 1
pub const ext_depth_clip_control_extension_name = "VK_EXT_depth_clip_control"
// PhysicalDeviceDepthClipControlFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDepthClipControlFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    depth_clip_control     Bool32
} 

// PipelineViewportDepthClipControlCreateInfoEXT extends VkPipelineViewportStateCreateInfo
pub struct PipelineViewportDepthClipControlCreateInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    negative_one_to_one    Bool32
} 



// VK_EXT_primitive_topology_list_restart is a preprocessor guard. Do not pass it to API calls.
const ext_primitive_topology_list_restart = 1
pub const ext_primitive_topology_list_restart_spec_version = 1
pub const ext_primitive_topology_list_restart_extension_name = "VK_EXT_primitive_topology_list_restart"
// PhysicalDevicePrimitiveTopologyListRestartFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePrimitiveTopologyListRestartFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    primitive_topology_list_restart Bool32
    primitive_topology_patch_list_restart Bool32
} 



// VK_FUCHSIA_external_memory is a preprocessor guard. Do not pass it to API calls.
const fuchsia_external_memory = 1
pub const fuchsia_external_memory_spec_version = 1
pub const fuchsia_external_memory_extension_name = "VK_CHSIA_external_memory"
// ImportMemoryZirconHandleInfoFUCHSIA extends VkMemoryAllocateInfo
pub struct ImportMemoryZirconHandleInfoFUCHSIA {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    handle_type                               ExternalMemoryHandleTypeFlagBits
    handle                                    voidptr
} 

pub struct MemoryZirconHandlePropertiesFUCHSIA {
mut:
    s_type                 StructureType
    p_next                 voidptr
    memory_type_bits       u32
} 

pub struct MemoryGetZirconHandleInfoFUCHSIA {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    memory                                    C.DeviceMemory
    handle_type                               ExternalMemoryHandleTypeFlagBits
} 

type VkGetMemoryZirconHandleFUCHSIA = fn (     C.Device,     &MemoryGetZirconHandleInfoFUCHSIA,     &voidptr) Result

pub fn get_memory_zircon_handle_fuchsia(
    device                                          C.Device,
    p_get_zircon_handle_info                        &MemoryGetZirconHandleInfoFUCHSIA,
    p_zircon_handle                                 &voidptr) Result {
      f := VkGetMemoryZirconHandleFUCHSIA((*loader_p).get_sym('vkGetMemoryZirconHandleFUCHSIA'
    ) or { 
        println("Couldn't load symbol for 'vkGetMemoryZirconHandleFUCHSIA': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_get_zircon_handle_info,
    p_zircon_handle)
}


type VkGetMemoryZirconHandlePropertiesFUCHSIA = fn (     C.Device,     ExternalMemoryHandleTypeFlagBits,     voidptr,     &MemoryZirconHandlePropertiesFUCHSIA) Result

pub fn get_memory_zircon_handle_properties_fuchsia(
    device                                          C.Device,
    handle_type                                     ExternalMemoryHandleTypeFlagBits,
    zircon_handle                                   voidptr,
    p_memory_zircon_handle_properties               &MemoryZirconHandlePropertiesFUCHSIA) Result {
      f := VkGetMemoryZirconHandlePropertiesFUCHSIA((*loader_p).get_sym('vkGetMemoryZirconHandlePropertiesFUCHSIA'
    ) or { 
        println("Couldn't load symbol for 'vkGetMemoryZirconHandlePropertiesFUCHSIA': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    handle_type,
    zircon_handle,
    p_memory_zircon_handle_properties)
}




// VK_FUCHSIA_external_semaphore is a preprocessor guard. Do not pass it to API calls.
const fuchsia_external_semaphore = 1
pub const fuchsia_external_semaphore_spec_version = 1
pub const fuchsia_external_semaphore_extension_name = "VK_CHSIA_external_semaphore"
pub struct ImportSemaphoreZirconHandleInfoFUCHSIA {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    semaphore                                    C.Semaphore
    flags                                        SemaphoreImportFlags
    handle_type                                  ExternalSemaphoreHandleTypeFlagBits
    zircon_handle                                voidptr
} 

pub struct SemaphoreGetZirconHandleInfoFUCHSIA {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    semaphore                                    C.Semaphore
    handle_type                                  ExternalSemaphoreHandleTypeFlagBits
} 

type VkImportSemaphoreZirconHandleFUCHSIA = fn (     C.Device,     &ImportSemaphoreZirconHandleInfoFUCHSIA) Result

pub fn import_semaphore_zircon_handle_fuchsia(
    device                                          C.Device,
    p_import_semaphore_zircon_handle_info           &ImportSemaphoreZirconHandleInfoFUCHSIA) Result {
      f := VkImportSemaphoreZirconHandleFUCHSIA((*loader_p).get_sym('vkImportSemaphoreZirconHandleFUCHSIA'
    ) or { 
        println("Couldn't load symbol for 'vkImportSemaphoreZirconHandleFUCHSIA': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_import_semaphore_zircon_handle_info)
}


type VkGetSemaphoreZirconHandleFUCHSIA = fn (     C.Device,     &SemaphoreGetZirconHandleInfoFUCHSIA,     &voidptr) Result

pub fn get_semaphore_zircon_handle_fuchsia(
    device                                          C.Device,
    p_get_zircon_handle_info                        &SemaphoreGetZirconHandleInfoFUCHSIA,
    p_zircon_handle                                 &voidptr) Result {
      f := VkGetSemaphoreZirconHandleFUCHSIA((*loader_p).get_sym('vkGetSemaphoreZirconHandleFUCHSIA'
    ) or { 
        println("Couldn't load symbol for 'vkGetSemaphoreZirconHandleFUCHSIA': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_get_zircon_handle_info,
    p_zircon_handle)
}




// VK_FUCHSIA_buffer_collection is a preprocessor guard. Do not pass it to API calls.
const fuchsia_buffer_collection = 1
pub type C.BufferCollectionFUCHSIA = voidptr
pub const fuchsia_buffer_collection_spec_version = 2
pub const fuchsia_buffer_collection_extension_name = "VK_CHSIA_buffer_collection"
pub type ImageFormatConstraintsFlagsFUCHSIA = u32

pub enum ImageConstraintsInfoFlagBitsFUCHSIA {
    image_constraints_info_cpu_read_rarely_fuchsia = int(0x00000001)
    image_constraints_info_cpu_read_often_fuchsia = int(0x00000002)
    image_constraints_info_cpu_write_rarely_fuchsia = int(0x00000004)
    image_constraints_info_cpu_write_often_fuchsia = int(0x00000008)
    image_constraints_info_protected_optional_fuchsia = int(0x00000010)
    image_constraints_info_flag_bits_max_enum_fuchsia = int(0x7FFFFFFF)
}

pub type ImageConstraintsInfoFlagsFUCHSIA = u32
pub struct BufferCollectionCreateInfoFUCHSIA {
mut:
    s_type                 StructureType
    p_next                 voidptr
    collection_token       voidptr
} 

// ImportMemoryBufferCollectionFUCHSIA extends VkMemoryAllocateInfo
pub struct ImportMemoryBufferCollectionFUCHSIA {
mut:
    s_type                           StructureType
    p_next                           voidptr
    collection                       C.BufferCollectionFUCHSIA
    index                            u32
} 

// BufferCollectionImageCreateInfoFUCHSIA extends VkImageCreateInfo
pub struct BufferCollectionImageCreateInfoFUCHSIA {
mut:
    s_type                           StructureType
    p_next                           voidptr
    collection                       C.BufferCollectionFUCHSIA
    index                            u32
} 

pub struct BufferCollectionConstraintsInfoFUCHSIA {
mut:
    s_type                 StructureType
    p_next                 voidptr
    min_buffer_count       u32
    max_buffer_count       u32
    min_buffer_count_for_camping u32
    min_buffer_count_for_dedicated_slack u32
    min_buffer_count_for_shared_slack u32
} 

pub struct BufferConstraintsInfoFUCHSIA {
mut:
    s_type                                          StructureType
    p_next                                          voidptr
    create_info                                     BufferCreateInfo
    required_format_features                        FormatFeatureFlags
    buffer_collection_constraints                   BufferCollectionConstraintsInfoFUCHSIA
} 

// BufferCollectionBufferCreateInfoFUCHSIA extends VkBufferCreateInfo
pub struct BufferCollectionBufferCreateInfoFUCHSIA {
mut:
    s_type                           StructureType
    p_next                           voidptr
    collection                       C.BufferCollectionFUCHSIA
    index                            u32
} 

pub struct SysmemColorSpaceFUCHSIA {
mut:
    s_type                 StructureType
    p_next                 voidptr
    color_space            u32
} 

pub struct BufferCollectionPropertiesFUCHSIA {
mut:
    s_type                               StructureType
    p_next                               voidptr
    memory_type_bits                     u32
    buffer_count                         u32
    create_info_index                    u32
    sysmem_pixel_format                  u64
    format_features                      FormatFeatureFlags
    sysmem_color_space_index             SysmemColorSpaceFUCHSIA
    sampler_ycbcr_conversion_components  ComponentMapping
    suggested_ycbcr_model                SamplerYcbcrModelConversion
    suggested_ycbcr_range                SamplerYcbcrRange
    suggested_x_chroma_offset            ChromaLocation
    suggested_y_chroma_offset            ChromaLocation
} 

pub struct ImageFormatConstraintsInfoFUCHSIA {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    image_create_info                           ImageCreateInfo
    required_format_features                    FormatFeatureFlags
    flags                                       ImageFormatConstraintsFlagsFUCHSIA
    sysmem_pixel_format                         u64
    color_space_count                           u32
    p_color_spaces                              &SysmemColorSpaceFUCHSIA
} 

pub struct ImageConstraintsInfoFUCHSIA {
mut:
    s_type                                            StructureType
    p_next                                            voidptr
    format_constraints_count                          u32
    p_format_constraints                              &ImageFormatConstraintsInfoFUCHSIA
    buffer_collection_constraints                     BufferCollectionConstraintsInfoFUCHSIA
    flags                                             ImageConstraintsInfoFlagsFUCHSIA
} 

type VkCreateBufferCollectionFUCHSIA = fn (     C.Device,     &BufferCollectionCreateInfoFUCHSIA,     &AllocationCallbacks,     &C.BufferCollectionFUCHSIA) Result

pub fn create_buffer_collection_fuchsia(
    device                                          C.Device,
    p_create_info                                   &BufferCollectionCreateInfoFUCHSIA,
    p_allocator                                     &AllocationCallbacks,
    p_collection                                    &C.BufferCollectionFUCHSIA) Result {
      f := VkCreateBufferCollectionFUCHSIA((*loader_p).get_sym('vkCreateBufferCollectionFUCHSIA'
    ) or { 
        println("Couldn't load symbol for 'vkCreateBufferCollectionFUCHSIA': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_collection)
}


type VkSetBufferCollectionImageConstraintsFUCHSIA = fn (     C.Device,     C.BufferCollectionFUCHSIA,     &ImageConstraintsInfoFUCHSIA) Result

pub fn set_buffer_collection_image_constraints_fuchsia(
    device                                          C.Device,
    collection                                      C.BufferCollectionFUCHSIA,
    p_image_constraints_info                        &ImageConstraintsInfoFUCHSIA) Result {
      f := VkSetBufferCollectionImageConstraintsFUCHSIA((*loader_p).get_sym('vkSetBufferCollectionImageConstraintsFUCHSIA'
    ) or { 
        println("Couldn't load symbol for 'vkSetBufferCollectionImageConstraintsFUCHSIA': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    collection,
    p_image_constraints_info)
}


type VkSetBufferCollectionBufferConstraintsFUCHSIA = fn (     C.Device,     C.BufferCollectionFUCHSIA,     &BufferConstraintsInfoFUCHSIA) Result

pub fn set_buffer_collection_buffer_constraints_fuchsia(
    device                                          C.Device,
    collection                                      C.BufferCollectionFUCHSIA,
    p_buffer_constraints_info                       &BufferConstraintsInfoFUCHSIA) Result {
      f := VkSetBufferCollectionBufferConstraintsFUCHSIA((*loader_p).get_sym('vkSetBufferCollectionBufferConstraintsFUCHSIA'
    ) or { 
        println("Couldn't load symbol for 'vkSetBufferCollectionBufferConstraintsFUCHSIA': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    collection,
    p_buffer_constraints_info)
}


type VkDestroyBufferCollectionFUCHSIA = fn (     C.Device,     C.BufferCollectionFUCHSIA,     &AllocationCallbacks) 

pub fn destroy_buffer_collection_fuchsia(
    device                                          C.Device,
    collection                                      C.BufferCollectionFUCHSIA,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyBufferCollectionFUCHSIA((*loader_p).get_sym('vkDestroyBufferCollectionFUCHSIA'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyBufferCollectionFUCHSIA': ${err}")
        return 
    })
    f(
    device,
    collection,
    p_allocator)
}


type VkGetBufferCollectionPropertiesFUCHSIA = fn (     C.Device,     C.BufferCollectionFUCHSIA,     &BufferCollectionPropertiesFUCHSIA) Result

pub fn get_buffer_collection_properties_fuchsia(
    device                                          C.Device,
    collection                                      C.BufferCollectionFUCHSIA,
    p_properties                                    &BufferCollectionPropertiesFUCHSIA) Result {
      f := VkGetBufferCollectionPropertiesFUCHSIA((*loader_p).get_sym('vkGetBufferCollectionPropertiesFUCHSIA'
    ) or { 
        println("Couldn't load symbol for 'vkGetBufferCollectionPropertiesFUCHSIA': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    collection,
    p_properties)
}




// VK_HUAWEI_subpass_shading is a preprocessor guard. Do not pass it to API calls.
const huawei_subpass_shading = 1
pub const huawei_subpass_shading_spec_version = 3
pub const huawei_subpass_shading_extension_name = "VK_HAWEI_subpass_shading"
// SubpassShadingPipelineCreateInfoHUAWEI extends VkComputePipelineCreateInfo
pub struct SubpassShadingPipelineCreateInfoHUAWEI {
mut:
    s_type                 StructureType
    p_next                 voidptr
    render_pass            C.RenderPass
    subpass                u32
} 

// PhysicalDeviceSubpassShadingFeaturesHUAWEI extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceSubpassShadingFeaturesHUAWEI {
mut:
    s_type                 StructureType
    p_next                 voidptr
    subpass_shading        Bool32
} 

// PhysicalDeviceSubpassShadingPropertiesHUAWEI extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceSubpassShadingPropertiesHUAWEI {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_subpass_shading_workgroup_size_aspect_ratio u32
} 

type VkGetDeviceSubpassShadingMaxWorkgroupSizeHUAWEI = fn (     C.Device,     C.RenderPass,     &Extent2D) Result

pub fn get_device_subpass_shading_max_workgroup_size_huawei(
    device                                          C.Device,
    renderpass                                      C.RenderPass,
    p_max_workgroup_size                            &Extent2D) Result {
      f := VkGetDeviceSubpassShadingMaxWorkgroupSizeHUAWEI((*loader_p).get_sym('vkGetDeviceSubpassShadingMaxWorkgroupSizeHUAWEI'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceSubpassShadingMaxWorkgroupSizeHUAWEI': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    renderpass,
    p_max_workgroup_size)
}


type VkCmdSubpassShadingHUAWEI = fn (     C.CommandBuffer) 

pub fn cmd_subpass_shading_huawei(
    command_buffer                                  C.CommandBuffer)  {
      f := VkCmdSubpassShadingHUAWEI((*loader_p).get_sym('vkCmdSubpassShadingHUAWEI'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSubpassShadingHUAWEI': ${err}")
        return 
    })
    f(
    command_buffer)
}




// VK_HUAWEI_invocation_mask is a preprocessor guard. Do not pass it to API calls.
const huawei_invocation_mask = 1
pub const huawei_invocation_mask_spec_version = 1
pub const huawei_invocation_mask_extension_name = "VK_HAWEI_invocation_mask"
// PhysicalDeviceInvocationMaskFeaturesHUAWEI extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceInvocationMaskFeaturesHUAWEI {
mut:
    s_type                 StructureType
    p_next                 voidptr
    invocation_mask        Bool32
} 

type VkCmdBindInvocationMaskHUAWEI = fn (     C.CommandBuffer,     C.ImageView,     ImageLayout) 

pub fn cmd_bind_invocation_mask_huawei(
    command_buffer                                  C.CommandBuffer,
    image_view                                      C.ImageView,
    image_layout                                    ImageLayout)  {
      f := VkCmdBindInvocationMaskHUAWEI((*loader_p).get_sym('vkCmdBindInvocationMaskHUAWEI'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindInvocationMaskHUAWEI': ${err}")
        return 
    })
    f(
    command_buffer,
    image_view,
    image_layout)
}




// VK_NV_external_memory_rdma is a preprocessor guard. Do not pass it to API calls.
const nv_external_memory_rdma = 1
pub type RemoteAddressNV = voidptr
pub const nv_external_memory_rdma_spec_version = 1
pub const nv_external_memory_rdma_extension_name = "VK_NV_external_memory_rdma"
pub struct MemoryGetRemoteAddressInfoNV {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    memory                                    C.DeviceMemory
    handle_type                               ExternalMemoryHandleTypeFlagBits
} 

// PhysicalDeviceExternalMemoryRDMAFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceExternalMemoryRDMAFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    external_memory_rdma   Bool32
} 

type VkGetMemoryRemoteAddressNV = fn (     C.Device,     &MemoryGetRemoteAddressInfoNV,     &RemoteAddressNV) Result

pub fn get_memory_remote_address_nv(
    device                                          C.Device,
    p_memory_get_remote_address_info                &MemoryGetRemoteAddressInfoNV,
    p_address                                       &RemoteAddressNV) Result {
      f := VkGetMemoryRemoteAddressNV((*loader_p).get_sym('vkGetMemoryRemoteAddressNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetMemoryRemoteAddressNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_memory_get_remote_address_info,
    p_address)
}




// VK_EXT_pipeline_properties is a preprocessor guard. Do not pass it to API calls.
const ext_pipeline_properties = 1
pub const ext_pipeline_properties_spec_version = 1
pub const ext_pipeline_properties_extension_name = "VK_EXT_pipeline_properties"
pub type PipelineInfoEXT = PipelineInfoKHR

pub struct PipelinePropertiesIdentifierEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pipeline_identifier    []u8
} 

// PhysicalDevicePipelinePropertiesFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePipelinePropertiesFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pipeline_properties_identifier Bool32
} 

type VkGetPipelinePropertiesEXT = fn (     C.Device,     &PipelineInfoEXT,     &BaseOutStructure) Result

pub fn get_pipeline_properties_ext(
    device                                          C.Device,
    p_pipeline_info                                 &PipelineInfoEXT,
    p_pipeline_properties                           &BaseOutStructure) Result {
      f := VkGetPipelinePropertiesEXT((*loader_p).get_sym('vkGetPipelinePropertiesEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetPipelinePropertiesEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_pipeline_info,
    p_pipeline_properties)
}




// VK_EXT_frame_boundary is a preprocessor guard. Do not pass it to API calls.
const ext_frame_boundary = 1
pub const ext_frame_boundary_spec_version   = 1
pub const ext_frame_boundary_extension_name = "VK_EXT_frame_boundary"

pub enum FrameBoundaryFlagBitsEXT {
    frame_boundary_frame_end_bit_ext = int(0x00000001)
    frame_boundary_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type FrameBoundaryFlagsEXT = u32
// PhysicalDeviceFrameBoundaryFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceFrameBoundaryFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    frame_boundary         Bool32
} 

// FrameBoundaryEXT extends VkSubmitInfo,VkSubmitInfo2,VkPresentInfoKHR,VkBindSparseInfo
pub struct FrameBoundaryEXT {
mut:
    s_type                         StructureType
    p_next                         voidptr
    flags                          FrameBoundaryFlagsEXT
    frame_id                       u64
    image_count                    u32
    p_images                       &C.Image
    buffer_count                   u32
    p_buffers                      &C.Buffer
    tag_name                       u64
    tag_size                       usize
    p_tag                          voidptr
} 



// VK_EXT_multisampled_render_to_single_sampled is a preprocessor guard. Do not pass it to API calls.
const ext_multisampled_render_to_single_sampled = 1
pub const ext_multisampled_render_to_single_sampled_spec_version = 1
pub const ext_multisampled_render_to_single_sampled_extension_name = "VK_EXT_multisampled_render_to_single_sampled"
// PhysicalDeviceMultisampledRenderToSingleSampledFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMultisampledRenderToSingleSampledFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    multisampled_render_to_single_sampled Bool32
} 

// SubpassResolvePerformanceQueryEXT extends VkFormatProperties2
pub struct SubpassResolvePerformanceQueryEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    optimal                Bool32
} 

// MultisampledRenderToSingleSampledInfoEXT extends VkSubpassDescription2,VkRenderingInfo
pub struct MultisampledRenderToSingleSampledInfoEXT {
mut:
    s_type                       StructureType
    p_next                       voidptr
    multisampled_render_to_single_sampled_enable Bool32
    rasterization_samples        SampleCountFlagBits
} 



// VK_EXT_extended_dynamic_state2 is a preprocessor guard. Do not pass it to API calls.
const ext_extended_dynamic_state2 = 1
pub const ext_extended_dynamic_state_2_spec_version = 1
pub const ext_extended_dynamic_state_2_extension_name = "VK_EXT_extended_dynamic_state2"
// PhysicalDeviceExtendedDynamicState2FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceExtendedDynamicState2FeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    extended_dynamic_state2 Bool32
    extended_dynamic_state2_logic_op Bool32
    extended_dynamic_state2_patch_control_points Bool32
} 

type VkCmdSetPatchControlPointsEXT = fn (     C.CommandBuffer,     u32) 

pub fn cmd_set_patch_control_points_ext(
    command_buffer                                  C.CommandBuffer,
    patch_control_points                            u32)  {
      f := VkCmdSetPatchControlPointsEXT((*loader_p).get_sym('vkCmdSetPatchControlPointsEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetPatchControlPointsEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    patch_control_points)
}


type VkCmdSetRasterizerDiscardEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_rasterizer_discard_enable_ext(
    command_buffer                                  C.CommandBuffer,
    rasterizer_discard_enable                       Bool32)  {
      f := VkCmdSetRasterizerDiscardEnableEXT((*loader_p).get_sym('vkCmdSetRasterizerDiscardEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetRasterizerDiscardEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    rasterizer_discard_enable)
}


type VkCmdSetDepthBiasEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_depth_bias_enable_ext(
    command_buffer                                  C.CommandBuffer,
    depth_bias_enable                               Bool32)  {
      f := VkCmdSetDepthBiasEnableEXT((*loader_p).get_sym('vkCmdSetDepthBiasEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthBiasEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_bias_enable)
}


type VkCmdSetLogicOpEXT = fn (     C.CommandBuffer,     LogicOp) 

pub fn cmd_set_logic_op_ext(
    command_buffer                                  C.CommandBuffer,
    logic_op                                        LogicOp)  {
      f := VkCmdSetLogicOpEXT((*loader_p).get_sym('vkCmdSetLogicOpEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetLogicOpEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    logic_op)
}


type VkCmdSetPrimitiveRestartEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_primitive_restart_enable_ext(
    command_buffer                                  C.CommandBuffer,
    primitive_restart_enable                        Bool32)  {
      f := VkCmdSetPrimitiveRestartEnableEXT((*loader_p).get_sym('vkCmdSetPrimitiveRestartEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetPrimitiveRestartEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    primitive_restart_enable)
}




// VK_QNX_screen_surface is a preprocessor guard. Do not pass it to API calls.
const qnx_screen_surface = 1
pub const qnx_screen_surface_spec_version   = 1
pub const qnx_screen_surface_extension_name = "VK_QNX_screen_surface"
pub type ScreenSurfaceCreateFlagsQNX = u32
pub struct ScreenSurfaceCreateInfoQNX {
mut:
    s_type                               StructureType
    p_next                               voidptr
    flags                                ScreenSurfaceCreateFlagsQNX
    context                              voidptr
    window                               voidptr
} 

type VkCreateScreenSurfaceQNX = fn (     C.Instance,     &ScreenSurfaceCreateInfoQNX,     &AllocationCallbacks,     &C.SurfaceKHR) Result

pub fn create_screen_surface_qnx(
    instance                                        C.Instance,
    p_create_info                                   &ScreenSurfaceCreateInfoQNX,
    p_allocator                                     &AllocationCallbacks,
    p_surface                                       &C.SurfaceKHR) Result {
      f := VkCreateScreenSurfaceQNX((*loader_p).get_sym('vkCreateScreenSurfaceQNX'
    ) or { 
        println("Couldn't load symbol for 'vkCreateScreenSurfaceQNX': ${err}")
        return Result.error_unknown
    })
    return f(
    instance,
    p_create_info,
    p_allocator,
    p_surface)
}


type VkGetPhysicalDeviceScreenPresentationSupportQNX = fn (     C.PhysicalDevice,     u32,     voidptr) Bool32

pub fn get_physical_device_screen_presentation_support_qnx(
    physical_device                                 C.PhysicalDevice,
    queue_family_index                              u32,
    window                                          voidptr) Bool32 {
      f := VkGetPhysicalDeviceScreenPresentationSupportQNX((*loader_p).get_sym("vkGetPhysicalDeviceScreenPresentationSupportQNX"
    ) or { 
        panic("Couldn't load symbol for 'vkGetPhysicalDeviceScreenPresentationSupportQNX': ${err}") })
    return f(
    physical_device,
    queue_family_index,
    window)
}




// VK_EXT_color_write_enable is a preprocessor guard. Do not pass it to API calls.
const ext_color_write_enable = 1
pub const ext_color_write_enable_spec_version = 1
pub const ext_color_write_enable_extension_name = "VK_EXT_color_write_enable"
// PhysicalDeviceColorWriteEnableFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceColorWriteEnableFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    color_write_enable     Bool32
} 

// PipelineColorWriteCreateInfoEXT extends VkPipelineColorBlendStateCreateInfo
pub struct PipelineColorWriteCreateInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    attachment_count       u32
    p_color_write_enables  &Bool32
} 

type VkCmdSetColorWriteEnableEXT = fn (     C.CommandBuffer,     u32,     &Bool32) 

pub fn cmd_set_color_write_enable_ext(
    command_buffer                                  C.CommandBuffer,
    attachment_count                                u32,
    p_color_write_enables                           &Bool32)  {
      f := VkCmdSetColorWriteEnableEXT((*loader_p).get_sym('vkCmdSetColorWriteEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetColorWriteEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    attachment_count,
    p_color_write_enables)
}




// VK_EXT_primitives_generated_query is a preprocessor guard. Do not pass it to API calls.
const ext_primitives_generated_query = 1
pub const ext_primitives_generated_query_spec_version = 1
pub const ext_primitives_generated_query_extension_name = "VK_EXT_primitives_generated_query"
// PhysicalDevicePrimitivesGeneratedQueryFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePrimitivesGeneratedQueryFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    primitives_generated_query Bool32
    primitives_generated_query_with_rasterizer_discard Bool32
    primitives_generated_query_with_non_zero_streams Bool32
} 



// VK_EXT_global_priority_query is a preprocessor guard. Do not pass it to API calls.
const ext_global_priority_query = 1
pub const ext_global_priority_query_spec_version = 1
pub const ext_global_priority_query_extension_name = "VK_EXT_global_priority_query"
pub const max_global_priority_size_ext      = max_global_priority_size_khr
pub type PhysicalDeviceGlobalPriorityQueryFeaturesEXT = PhysicalDeviceGlobalPriorityQueryFeaturesKHR

pub type QueueFamilyGlobalPriorityPropertiesEXT = QueueFamilyGlobalPriorityPropertiesKHR



// VK_EXT_image_view_min_lod is a preprocessor guard. Do not pass it to API calls.
const ext_image_view_min_lod = 1
pub const ext_image_view_min_lod_spec_version = 1
pub const ext_image_view_min_lod_extension_name = "VK_EXT_image_view_min_lod"
// PhysicalDeviceImageViewMinLodFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceImageViewMinLodFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    min_lod                Bool32
} 

// ImageViewMinLodCreateInfoEXT extends VkImageViewCreateInfo
pub struct ImageViewMinLodCreateInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    min_lod                f32
} 



// VK_EXT_multi_draw is a preprocessor guard. Do not pass it to API calls.
const ext_multi_draw = 1
pub const ext_multi_draw_spec_version       = 1
pub const ext_multi_draw_extension_name     = "VK_EXT_multi_draw"
// PhysicalDeviceMultiDrawFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMultiDrawFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    multi_draw             Bool32
} 

// PhysicalDeviceMultiDrawPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceMultiDrawPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_multi_draw_count   u32
} 

pub struct MultiDrawInfoEXT {
mut:
    first_vertex    u32
    vertex_count    u32
} 

pub struct MultiDrawIndexedInfoEXT {
mut:
    first_index     u32
    index_count     u32
    vertex_offset   i32
} 

type VkCmdDrawMultiEXT = fn (     C.CommandBuffer,     u32,     &MultiDrawInfoEXT,     u32,     u32,     u32) 

pub fn cmd_draw_multi_ext(
    command_buffer                                  C.CommandBuffer,
    draw_count                                      u32,
    p_vertex_info                                   &MultiDrawInfoEXT,
    instance_count                                  u32,
    first_instance                                  u32,
    stride                                          u32)  {
      f := VkCmdDrawMultiEXT((*loader_p).get_sym('vkCmdDrawMultiEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawMultiEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    draw_count,
    p_vertex_info,
    instance_count,
    first_instance,
    stride)
}


type VkCmdDrawMultiIndexedEXT = fn (     C.CommandBuffer,     u32,     &MultiDrawIndexedInfoEXT,     u32,     u32,     u32,     &i32) 

pub fn cmd_draw_multi_indexed_ext(
    command_buffer                                  C.CommandBuffer,
    draw_count                                      u32,
    p_index_info                                    &MultiDrawIndexedInfoEXT,
    instance_count                                  u32,
    first_instance                                  u32,
    stride                                          u32,
    p_vertex_offset                                 &i32)  {
      f := VkCmdDrawMultiIndexedEXT((*loader_p).get_sym('vkCmdDrawMultiIndexedEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawMultiIndexedEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    draw_count,
    p_index_info,
    instance_count,
    first_instance,
    stride,
    p_vertex_offset)
}




// VK_EXT_image_2d_view_of_3d is a preprocessor guard. Do not pass it to API calls.
const ext_image_2d_view_of_3d = 1
pub const ext_image_2d_view_of_3d_spec_version = 1
pub const ext_image_2d_view_of_3d_extension_name = "VK_EXT_image_2d_view_of_3d"
// PhysicalDeviceImage2DViewOf3DFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceImage2DViewOf3DFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image2_d_view_of3_d    Bool32
    sampler2_d_view_of3_d  Bool32
} 



// VK_EXT_shader_tile_image is a preprocessor guard. Do not pass it to API calls.
const ext_shader_tile_image = 1
pub const ext_shader_tile_image_spec_version = 1
pub const ext_shader_tile_image_extension_name = "VK_EXT_shader_tile_image"
// PhysicalDeviceShaderTileImageFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderTileImageFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_tile_image_color_read_access Bool32
    shader_tile_image_depth_read_access Bool32
    shader_tile_image_stencil_read_access Bool32
} 

// PhysicalDeviceShaderTileImagePropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceShaderTileImagePropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_tile_image_coherent_read_accelerated Bool32
    shader_tile_image_read_sample_from_pixel_rate_invocation Bool32
    shader_tile_image_read_from_helper_invocation Bool32
} 



// VK_EXT_opacity_micromap is a preprocessor guard. Do not pass it to API calls.
const ext_opacity_micromap = 1
pub type C.MicromapEXT = voidptr
pub const ext_opacity_micromap_spec_version = 2
pub const ext_opacity_micromap_extension_name = "VK_EXT_opacity_micromap"

pub enum MicromapTypeEXT {
    micromap_type_opacity_micromap_ext = int(0)
    micromap_type_max_enum_ext = int(0x7FFFFFFF)
}


pub enum BuildMicromapModeEXT {
    build_micromap_mode_build_ext = int(0)
    build_micromap_mode_max_enum_ext = int(0x7FFFFFFF)
}


pub enum CopyMicromapModeEXT {
    copy_micromap_mode_clone_ext = int(0)
    copy_micromap_mode_serialize_ext = int(1)
    copy_micromap_mode_deserialize_ext = int(2)
    copy_micromap_mode_compact_ext = int(3)
    copy_micromap_mode_max_enum_ext = int(0x7FFFFFFF)
}


pub enum OpacityMicromapFormatEXT {
    opacity_micromap_format_2_state_ext = int(1)
    opacity_micromap_format_4_state_ext = int(2)
    opacity_micromap_format_max_enum_ext = int(0x7FFFFFFF)
}


pub enum OpacityMicromapSpecialIndexEXT {
    opacity_micromap_special_index_fully_transparent_ext = int(-1)
    opacity_micromap_special_index_fully_opaque_ext = int(-2)
    opacity_micromap_special_index_fully_unknown_transparent_ext = int(-3)
    opacity_micromap_special_index_fully_unknown_opaque_ext = int(-4)
    opacity_micromap_special_index_max_enum_ext = int(0x7FFFFFFF)
}


pub enum AccelerationStructureCompatibilityKHR {
    acceleration_structure_compatibility_compatible_khr = int(0)
    acceleration_structure_compatibility_incompatible_khr = int(1)
    acceleration_structure_compatibility_max_enum_khr = int(0x7FFFFFFF)
}


pub enum AccelerationStructureBuildTypeKHR {
    acceleration_structure_build_type_host_khr = int(0)
    acceleration_structure_build_type_device_khr = int(1)
    acceleration_structure_build_type_host_or_device_khr = int(2)
    acceleration_structure_build_type_max_enum_khr = int(0x7FFFFFFF)
}


pub enum BuildMicromapFlagBitsEXT {
    build_micromap_prefer_fast_trace_bit_ext = int(0x00000001)
    build_micromap_prefer_fast_build_bit_ext = int(0x00000002)
    build_micromap_allow_compaction_bit_ext = int(0x00000004)
    build_micromap_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type BuildMicromapFlagsEXT = u32

pub enum MicromapCreateFlagBitsEXT {
    micromap_create_device_address_capture_replay_bit_ext = int(0x00000001)
    micromap_create_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type MicromapCreateFlagsEXT = u32
pub struct MicromapUsageEXT {
mut:
    count           u32
    subdivision_level u32
    format          u32
} 

pub union DeviceOrHostAddressKHR {
mut:
    device_address         DeviceAddress
    host_address           voidptr
} 

pub struct MicromapBuildInfoEXT {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    vktype                                  MicromapTypeEXT
    flags                                   BuildMicromapFlagsEXT
    mode                                    BuildMicromapModeEXT
    dst_micromap                            C.MicromapEXT
    usage_counts_count                      u32
    p_usage_counts                          &MicromapUsageEXT
    pp_usage_counts                         &MicromapUsageEXT
    data                                    DeviceOrHostAddressConstKHR
    scratch_data                            DeviceOrHostAddressKHR
    triangle_array                          DeviceOrHostAddressConstKHR
    triangle_array_stride                   DeviceSize
} 

pub struct MicromapCreateInfoEXT {
mut:
    s_type                          StructureType
    p_next                          voidptr
    create_flags                    MicromapCreateFlagsEXT
    buffer                          C.Buffer
    offset                          DeviceSize
    size                            DeviceSize
    vktype                          MicromapTypeEXT
    device_address                  DeviceAddress
} 

// PhysicalDeviceOpacityMicromapFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceOpacityMicromapFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    micromap               Bool32
    micromap_capture_replay Bool32
    micromap_host_commands Bool32
} 

// PhysicalDeviceOpacityMicromapPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceOpacityMicromapPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_opacity2_state_subdivision_level u32
    max_opacity4_state_subdivision_level u32
} 

pub struct MicromapVersionInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    p_version_data         &u8
} 

pub struct CopyMicromapToMemoryInfoEXT {
mut:
    s_type                          StructureType
    p_next                          voidptr
    src                             C.MicromapEXT
    dst                             DeviceOrHostAddressKHR
    mode                            CopyMicromapModeEXT
} 

pub struct CopyMemoryToMicromapInfoEXT {
mut:
    s_type                               StructureType
    p_next                               voidptr
    src                                  DeviceOrHostAddressConstKHR
    dst                                  C.MicromapEXT
    mode                                 CopyMicromapModeEXT
} 

pub struct CopyMicromapInfoEXT {
mut:
    s_type                       StructureType
    p_next                       voidptr
    src                          C.MicromapEXT
    dst                          C.MicromapEXT
    mode                         CopyMicromapModeEXT
} 

pub struct MicromapBuildSizesInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    micromap_size          DeviceSize
    build_scratch_size     DeviceSize
    discardable            Bool32
} 

// AccelerationStructureTrianglesOpacityMicromapEXT extends VkAccelerationStructureGeometryTrianglesDataKHR
pub struct AccelerationStructureTrianglesOpacityMicromapEXT {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    index_type                              IndexType
    index_buffer                            DeviceOrHostAddressConstKHR
    index_stride                            DeviceSize
    base_triangle                           u32
    usage_counts_count                      u32
    p_usage_counts                          &MicromapUsageEXT
    pp_usage_counts                         &MicromapUsageEXT
    micromap                                C.MicromapEXT
} 

pub struct MicromapTriangleEXT {
mut:
    data_offset     u32
    subdivision_level u16
    format          u16
} 

type VkCreateMicromapEXT = fn (     C.Device,     &MicromapCreateInfoEXT,     &AllocationCallbacks,     &C.MicromapEXT) Result

pub fn create_micromap_ext(
    device                                          C.Device,
    p_create_info                                   &MicromapCreateInfoEXT,
    p_allocator                                     &AllocationCallbacks,
    p_micromap                                      &C.MicromapEXT) Result {
      f := VkCreateMicromapEXT((*loader_p).get_sym('vkCreateMicromapEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCreateMicromapEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_micromap)
}


type VkDestroyMicromapEXT = fn (     C.Device,     C.MicromapEXT,     &AllocationCallbacks) 

pub fn destroy_micromap_ext(
    device                                          C.Device,
    micromap                                        C.MicromapEXT,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyMicromapEXT((*loader_p).get_sym('vkDestroyMicromapEXT'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyMicromapEXT': ${err}")
        return 
    })
    f(
    device,
    micromap,
    p_allocator)
}


type VkCmdBuildMicromapsEXT = fn (     C.CommandBuffer,     u32,     &MicromapBuildInfoEXT) 

pub fn cmd_build_micromaps_ext(
    command_buffer                                  C.CommandBuffer,
    info_count                                      u32,
    p_infos                                         &MicromapBuildInfoEXT)  {
      f := VkCmdBuildMicromapsEXT((*loader_p).get_sym('vkCmdBuildMicromapsEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBuildMicromapsEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    info_count,
    p_infos)
}


type VkBuildMicromapsEXT = fn (     C.Device,     C.DeferredOperationKHR,     u32,     &MicromapBuildInfoEXT) Result

pub fn build_micromaps_ext(
    device                                          C.Device,
    deferred_operation                              C.DeferredOperationKHR,
    info_count                                      u32,
    p_infos                                         &MicromapBuildInfoEXT) Result {
      f := VkBuildMicromapsEXT((*loader_p).get_sym('vkBuildMicromapsEXT'
    ) or { 
        println("Couldn't load symbol for 'vkBuildMicromapsEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    deferred_operation,
    info_count,
    p_infos)
}


type VkCopyMicromapEXT = fn (     C.Device,     C.DeferredOperationKHR,     &CopyMicromapInfoEXT) Result

pub fn copy_micromap_ext(
    device                                          C.Device,
    deferred_operation                              C.DeferredOperationKHR,
    p_info                                          &CopyMicromapInfoEXT) Result {
      f := VkCopyMicromapEXT((*loader_p).get_sym('vkCopyMicromapEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCopyMicromapEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    deferred_operation,
    p_info)
}


type VkCopyMicromapToMemoryEXT = fn (     C.Device,     C.DeferredOperationKHR,     &CopyMicromapToMemoryInfoEXT) Result

pub fn copy_micromap_to_memory_ext(
    device                                          C.Device,
    deferred_operation                              C.DeferredOperationKHR,
    p_info                                          &CopyMicromapToMemoryInfoEXT) Result {
      f := VkCopyMicromapToMemoryEXT((*loader_p).get_sym('vkCopyMicromapToMemoryEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCopyMicromapToMemoryEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    deferred_operation,
    p_info)
}


type VkCopyMemoryToMicromapEXT = fn (     C.Device,     C.DeferredOperationKHR,     &CopyMemoryToMicromapInfoEXT) Result

pub fn copy_memory_to_micromap_ext(
    device                                          C.Device,
    deferred_operation                              C.DeferredOperationKHR,
    p_info                                          &CopyMemoryToMicromapInfoEXT) Result {
      f := VkCopyMemoryToMicromapEXT((*loader_p).get_sym('vkCopyMemoryToMicromapEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCopyMemoryToMicromapEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    deferred_operation,
    p_info)
}


type VkWriteMicromapsPropertiesEXT = fn (     C.Device,     u32,     &C.MicromapEXT,     QueryType,     usize,     voidptr,     usize) Result

pub fn write_micromaps_properties_ext(
    device                                          C.Device,
    micromap_count                                  u32,
    p_micromaps                                     &C.MicromapEXT,
    query_type                                      QueryType,
    data_size                                       usize,
    p_data                                          voidptr,
    stride                                          usize) Result {
      f := VkWriteMicromapsPropertiesEXT((*loader_p).get_sym('vkWriteMicromapsPropertiesEXT'
    ) or { 
        println("Couldn't load symbol for 'vkWriteMicromapsPropertiesEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    micromap_count,
    p_micromaps,
    query_type,
    data_size,
    p_data,
    stride)
}


type VkCmdCopyMicromapEXT = fn (     C.CommandBuffer,     &CopyMicromapInfoEXT) 

pub fn cmd_copy_micromap_ext(
    command_buffer                                  C.CommandBuffer,
    p_info                                          &CopyMicromapInfoEXT)  {
      f := VkCmdCopyMicromapEXT((*loader_p).get_sym('vkCmdCopyMicromapEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyMicromapEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    p_info)
}


type VkCmdCopyMicromapToMemoryEXT = fn (     C.CommandBuffer,     &CopyMicromapToMemoryInfoEXT) 

pub fn cmd_copy_micromap_to_memory_ext(
    command_buffer                                  C.CommandBuffer,
    p_info                                          &CopyMicromapToMemoryInfoEXT)  {
      f := VkCmdCopyMicromapToMemoryEXT((*loader_p).get_sym('vkCmdCopyMicromapToMemoryEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyMicromapToMemoryEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    p_info)
}


type VkCmdCopyMemoryToMicromapEXT = fn (     C.CommandBuffer,     &CopyMemoryToMicromapInfoEXT) 

pub fn cmd_copy_memory_to_micromap_ext(
    command_buffer                                  C.CommandBuffer,
    p_info                                          &CopyMemoryToMicromapInfoEXT)  {
      f := VkCmdCopyMemoryToMicromapEXT((*loader_p).get_sym('vkCmdCopyMemoryToMicromapEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyMemoryToMicromapEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    p_info)
}


type VkCmdWriteMicromapsPropertiesEXT = fn (     C.CommandBuffer,     u32,     &C.MicromapEXT,     QueryType,     C.QueryPool,     u32) 

pub fn cmd_write_micromaps_properties_ext(
    command_buffer                                  C.CommandBuffer,
    micromap_count                                  u32,
    p_micromaps                                     &C.MicromapEXT,
    query_type                                      QueryType,
    query_pool                                      C.QueryPool,
    first_query                                     u32)  {
      f := VkCmdWriteMicromapsPropertiesEXT((*loader_p).get_sym('vkCmdWriteMicromapsPropertiesEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdWriteMicromapsPropertiesEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    micromap_count,
    p_micromaps,
    query_type,
    query_pool,
    first_query)
}


type VkGetDeviceMicromapCompatibilityEXT = fn (     C.Device,     &MicromapVersionInfoEXT,     &AccelerationStructureCompatibilityKHR) 

pub fn get_device_micromap_compatibility_ext(
    device                                          C.Device,
    p_version_info                                  &MicromapVersionInfoEXT,
    p_compatibility                                 &AccelerationStructureCompatibilityKHR)  {
      f := VkGetDeviceMicromapCompatibilityEXT((*loader_p).get_sym('vkGetDeviceMicromapCompatibilityEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceMicromapCompatibilityEXT': ${err}")
        return 
    })
    f(
    device,
    p_version_info,
    p_compatibility)
}


type VkGetMicromapBuildSizesEXT = fn (     C.Device,     AccelerationStructureBuildTypeKHR,     &MicromapBuildInfoEXT,     &MicromapBuildSizesInfoEXT) 

pub fn get_micromap_build_sizes_ext(
    device                                          C.Device,
    build_type                                      AccelerationStructureBuildTypeKHR,
    p_build_info                                    &MicromapBuildInfoEXT,
    p_size_info                                     &MicromapBuildSizesInfoEXT)  {
      f := VkGetMicromapBuildSizesEXT((*loader_p).get_sym('vkGetMicromapBuildSizesEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetMicromapBuildSizesEXT': ${err}")
        return 
    })
    f(
    device,
    build_type,
    p_build_info,
    p_size_info)
}




// VK_NV_displacement_micromap is a preprocessor guard. Do not pass it to API calls.
const nv_displacement_micromap = 1
pub const nv_displacement_micromap_spec_version = 2
pub const nv_displacement_micromap_extension_name = "VK_NV_displacement_micromap"

pub enum DisplacementMicromapFormatNV {
    displacement_micromap_format_64_triangles_64_bytes_nv = int(1)
    displacement_micromap_format_256_triangles_128_bytes_nv = int(2)
    displacement_micromap_format_1024_triangles_128_bytes_nv = int(3)
    displacement_micromap_format_max_enum_nv = int(0x7FFFFFFF)
}

// PhysicalDeviceDisplacementMicromapFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDisplacementMicromapFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    displacement_micromap  Bool32
} 

// PhysicalDeviceDisplacementMicromapPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceDisplacementMicromapPropertiesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_displacement_micromap_subdivision_level u32
} 

// AccelerationStructureTrianglesDisplacementMicromapNV extends VkAccelerationStructureGeometryTrianglesDataKHR
pub struct AccelerationStructureTrianglesDisplacementMicromapNV {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    displacement_bias_and_scale_format      Format
    displacement_vector_format              Format
    displacement_bias_and_scale_buffer      DeviceOrHostAddressConstKHR
    displacement_bias_and_scale_stride      DeviceSize
    displacement_vector_buffer              DeviceOrHostAddressConstKHR
    displacement_vector_stride              DeviceSize
    displaced_micromap_primitive_flags      DeviceOrHostAddressConstKHR
    displaced_micromap_primitive_flags_stride DeviceSize
    index_type                              IndexType
    index_buffer                            DeviceOrHostAddressConstKHR
    index_stride                            DeviceSize
    base_triangle                           u32
    usage_counts_count                      u32
    p_usage_counts                          &MicromapUsageEXT
    pp_usage_counts                         &MicromapUsageEXT
    micromap                                C.MicromapEXT
} 



// VK_EXT_load_store_op_none is a preprocessor guard. Do not pass it to API calls.
const ext_load_store_op_none = 1
pub const ext_load_store_op_none_spec_version = 1
pub const ext_load_store_op_none_extension_name = "VK_EXT_load_store_op_none"


// VK_HUAWEI_cluster_culling_shader is a preprocessor guard. Do not pass it to API calls.
const huawei_cluster_culling_shader = 1
pub const huawei_cluster_culling_shader_spec_version = 3
pub const huawei_cluster_culling_shader_extension_name = "VK_HAWEI_cluster_culling_shader"
// PhysicalDeviceClusterCullingShaderFeaturesHUAWEI extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceClusterCullingShaderFeaturesHUAWEI {
mut:
    s_type                 StructureType
    p_next                 voidptr
    clusterculling_shader  Bool32
    multiview_cluster_culling_shader Bool32
} 

// PhysicalDeviceClusterCullingShaderPropertiesHUAWEI extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceClusterCullingShaderPropertiesHUAWEI {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_work_group_count   []u32
    max_work_group_size    []u32
    max_output_cluster_count u32
    indirect_buffer_offset_alignment DeviceSize
} 

// PhysicalDeviceClusterCullingShaderVrsFeaturesHUAWEI extends VkPhysicalDeviceClusterCullingShaderFeaturesHUAWEI
pub struct PhysicalDeviceClusterCullingShaderVrsFeaturesHUAWEI {
mut:
    s_type                 StructureType
    p_next                 voidptr
    cluster_shading_rate   Bool32
} 

type VkCmdDrawClusterHUAWEI = fn (     C.CommandBuffer,     u32,     u32,     u32) 

pub fn cmd_draw_cluster_huawei(
    command_buffer                                  C.CommandBuffer,
    group_count_x                                   u32,
    group_count_y                                   u32,
    group_count_z                                   u32)  {
      f := VkCmdDrawClusterHUAWEI((*loader_p).get_sym('vkCmdDrawClusterHUAWEI'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawClusterHUAWEI': ${err}")
        return 
    })
    f(
    command_buffer,
    group_count_x,
    group_count_y,
    group_count_z)
}


type VkCmdDrawClusterIndirectHUAWEI = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize) 

pub fn cmd_draw_cluster_indirect_huawei(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize)  {
      f := VkCmdDrawClusterIndirectHUAWEI((*loader_p).get_sym('vkCmdDrawClusterIndirectHUAWEI'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawClusterIndirectHUAWEI': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset)
}




// VK_EXT_border_color_swizzle is a preprocessor guard. Do not pass it to API calls.
const ext_border_color_swizzle = 1
pub const ext_border_color_swizzle_spec_version = 1
pub const ext_border_color_swizzle_extension_name = "VK_EXT_border_color_swizzle"
// PhysicalDeviceBorderColorSwizzleFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceBorderColorSwizzleFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    border_color_swizzle   Bool32
    border_color_swizzle_from_image Bool32
} 

// SamplerBorderColorComponentMappingCreateInfoEXT extends VkSamplerCreateInfo
pub struct SamplerBorderColorComponentMappingCreateInfoEXT {
mut:
    s_type                    StructureType
    p_next                    voidptr
    components                ComponentMapping
    srgb                      Bool32
} 



// VK_EXT_pageable_device_local_memory is a preprocessor guard. Do not pass it to API calls.
const ext_pageable_device_local_memory = 1
pub const ext_pageable_device_local_memory_spec_version = 1
pub const ext_pageable_device_local_memory_extension_name = "VK_EXT_pageable_device_local_memory"
// PhysicalDevicePageableDeviceLocalMemoryFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePageableDeviceLocalMemoryFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pageable_device_local_memory Bool32
} 

type VkSetDeviceMemoryPriorityEXT = fn (     C.Device,     C.DeviceMemory,     f32) 

pub fn set_device_memory_priority_ext(
    device                                          C.Device,
    memory                                          C.DeviceMemory,
    priority                                        f32)  {
      f := VkSetDeviceMemoryPriorityEXT((*loader_p).get_sym('vkSetDeviceMemoryPriorityEXT'
    ) or { 
        println("Couldn't load symbol for 'vkSetDeviceMemoryPriorityEXT': ${err}")
        return 
    })
    f(
    device,
    memory,
    priority)
}




// VK_ARM_shader_core_properties is a preprocessor guard. Do not pass it to API calls.
const arm_shader_core_properties = 1
pub const arm_shader_core_properties_spec_version = 1
pub const arm_shader_core_properties_extension_name = "VK_ARM_shader_core_properties"
// PhysicalDeviceShaderCorePropertiesARM extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceShaderCorePropertiesARM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pixel_rate             u32
    texel_rate             u32
    fma_rate               u32
} 



// VK_ARM_scheduling_controls is a preprocessor guard. Do not pass it to API calls.
const arm_scheduling_controls = 1
pub const arm_scheduling_controls_spec_version = 1
pub const arm_scheduling_controls_extension_name = "VK_ARM_scheduling_controls"
pub type PhysicalDeviceSchedulingControlsFlagsARM = u64

pub enum PhysicalDeviceSchedulingControlsFlagBitsARM {
    physical_device_scheduling_controls_shader_core_count_arm = int(0x00000001)
    physical_device_scheduling_controls_flag_bits_max_enum_arm = int(0x7FFFFFFF)
}

// DeviceQueueShaderCoreControlCreateInfoARM extends VkDeviceQueueCreateInfo,VkDeviceCreateInfo
pub struct DeviceQueueShaderCoreControlCreateInfoARM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_core_count      u32
} 

// PhysicalDeviceSchedulingControlsFeaturesARM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceSchedulingControlsFeaturesARM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    scheduling_controls    Bool32
} 

// PhysicalDeviceSchedulingControlsPropertiesARM extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceSchedulingControlsPropertiesARM {
mut:
    s_type                                            StructureType
    p_next                                            voidptr
    scheduling_controls_flags                         PhysicalDeviceSchedulingControlsFlagsARM
} 



// VK_EXT_image_sliced_view_of_3d is a preprocessor guard. Do not pass it to API calls.
const ext_image_sliced_view_of_3d = 1
pub const ext_image_sliced_view_of_3d_spec_version = 1
pub const ext_image_sliced_view_of_3d_extension_name = "VK_EXT_image_sliced_view_of_3d"
pub const remaining_3d_slices_ext           = ~u32(0)
// PhysicalDeviceImageSlicedViewOf3DFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceImageSlicedViewOf3DFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image_sliced_view_of3_d Bool32
} 

// ImageViewSlicedCreateInfoEXT extends VkImageViewCreateInfo
pub struct ImageViewSlicedCreateInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    slice_offset           u32
    slice_count            u32
} 



// VK_VALVE_descriptor_set_host_mapping is a preprocessor guard. Do not pass it to API calls.
const valve_descriptor_set_host_mapping = 1
pub const valve_descriptor_set_host_mapping_spec_version = 1
pub const valve_descriptor_set_host_mapping_extension_name = "VK_VAVE_descriptor_set_host_mapping"
// PhysicalDeviceDescriptorSetHostMappingFeaturesVALVE extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDescriptorSetHostMappingFeaturesVALVE {
mut:
    s_type                 StructureType
    p_next                 voidptr
    descriptor_set_host_mapping Bool32
} 

pub struct DescriptorSetBindingReferenceVALVE {
mut:
    s_type                       StructureType
    p_next                       voidptr
    descriptor_set_layout        C.DescriptorSetLayout
    binding                      u32
} 

pub struct DescriptorSetLayoutHostMappingInfoVALVE {
mut:
    s_type                 StructureType
    p_next                 voidptr
    descriptor_offset      usize
    descriptor_size        u32
} 

type VkGetDescriptorSetLayoutHostMappingInfoVALVE = fn (     C.Device,     &DescriptorSetBindingReferenceVALVE,     &DescriptorSetLayoutHostMappingInfoVALVE) 

pub fn get_descriptor_set_layout_host_mapping_info_valve(
    device                                          C.Device,
    p_binding_reference                             &DescriptorSetBindingReferenceVALVE,
    p_host_mapping                                  &DescriptorSetLayoutHostMappingInfoVALVE)  {
      f := VkGetDescriptorSetLayoutHostMappingInfoVALVE((*loader_p).get_sym('vkGetDescriptorSetLayoutHostMappingInfoVALVE'
    ) or { 
        println("Couldn't load symbol for 'vkGetDescriptorSetLayoutHostMappingInfoVALVE': ${err}")
        return 
    })
    f(
    device,
    p_binding_reference,
    p_host_mapping)
}


type VkGetDescriptorSetHostMappingVALVE = fn (     C.Device,     C.DescriptorSet,     &voidptr) 

pub fn get_descriptor_set_host_mapping_valve(
    device                                          C.Device,
    descriptor_set                                  C.DescriptorSet,
    pp_data                                         &voidptr)  {
      f := VkGetDescriptorSetHostMappingVALVE((*loader_p).get_sym('vkGetDescriptorSetHostMappingVALVE'
    ) or { 
        println("Couldn't load symbol for 'vkGetDescriptorSetHostMappingVALVE': ${err}")
        return 
    })
    f(
    device,
    descriptor_set,
    pp_data)
}




// VK_EXT_depth_clamp_zero_one is a preprocessor guard. Do not pass it to API calls.
const ext_depth_clamp_zero_one = 1
pub const ext_depth_clamp_zero_one_spec_version = 1
pub const ext_depth_clamp_zero_one_extension_name = "VK_EXT_depth_clamp_zero_one"
// PhysicalDeviceDepthClampZeroOneFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDepthClampZeroOneFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    depth_clamp_zero_one   Bool32
} 



// VK_EXT_non_seamless_cube_map is a preprocessor guard. Do not pass it to API calls.
const ext_non_seamless_cube_map = 1
pub const ext_non_seamless_cube_map_spec_version = 1
pub const ext_non_seamless_cube_map_extension_name = "VK_EXT_non_seamless_cube_map"
// PhysicalDeviceNonSeamlessCubeMapFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceNonSeamlessCubeMapFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    non_seamless_cube_map  Bool32
} 



// VK_ARM_render_pass_striped is a preprocessor guard. Do not pass it to API calls.
const arm_render_pass_striped = 1
pub const arm_render_pass_striped_spec_version = 1
pub const arm_render_pass_striped_extension_name = "VK_ARM_render_pass_striped"
// PhysicalDeviceRenderPassStripedFeaturesARM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRenderPassStripedFeaturesARM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    render_pass_striped    Bool32
} 

// PhysicalDeviceRenderPassStripedPropertiesARM extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceRenderPassStripedPropertiesARM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    render_pass_stripe_granularity Extent2D
    max_render_pass_stripes u32
} 

pub struct RenderPassStripeInfoARM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    stripe_area            Rect2D
} 

// RenderPassStripeBeginInfoARM extends VkRenderingInfo,VkRenderPassBeginInfo
pub struct RenderPassStripeBeginInfoARM {
mut:
    s_type                            StructureType
    p_next                            voidptr
    stripe_info_count                 u32
    p_stripe_infos                    &RenderPassStripeInfoARM
} 

// RenderPassStripeSubmitInfoARM extends VkCommandBufferSubmitInfo
pub struct RenderPassStripeSubmitInfoARM {
mut:
    s_type                              StructureType
    p_next                              voidptr
    stripe_semaphore_info_count         u32
    p_stripe_semaphore_infos            &SemaphoreSubmitInfo
} 



// VK_QCOM_fragment_density_map_offset is a preprocessor guard. Do not pass it to API calls.
const qcom_fragment_density_map_offset = 1
pub const qcom_fragment_density_map_offset_spec_version = 1
pub const qcom_fragment_density_map_offset_extension_name = "VK_QCOM_fragment_density_map_offset"
// PhysicalDeviceFragmentDensityMapOffsetFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceFragmentDensityMapOffsetFeaturesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    fragment_density_map_offset Bool32
} 

// PhysicalDeviceFragmentDensityMapOffsetPropertiesQCOM extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceFragmentDensityMapOffsetPropertiesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    fragment_density_offset_granularity Extent2D
} 

// SubpassFragmentDensityMapOffsetEndInfoQCOM extends VkSubpassEndInfo
pub struct SubpassFragmentDensityMapOffsetEndInfoQCOM {
mut:
    s_type                   StructureType
    p_next                   voidptr
    fragment_density_offset_count u32
    p_fragment_density_offsets &Offset2D
} 



// VK_NV_copy_memory_indirect is a preprocessor guard. Do not pass it to API calls.
const nv_copy_memory_indirect = 1
pub const nv_copy_memory_indirect_spec_version = 1
pub const nv_copy_memory_indirect_extension_name = "VK_NV_copy_memory_indirect"
pub struct CopyMemoryIndirectCommandNV {
mut:
    src_address            DeviceAddress
    dst_address            DeviceAddress
    size                   DeviceSize
} 

pub struct CopyMemoryToImageIndirectCommandNV {
mut:
    src_address                     DeviceAddress
    buffer_row_length               u32
    buffer_image_height             u32
    image_subresource               ImageSubresourceLayers
    image_offset                    Offset3D
    image_extent                    Extent3D
} 

// PhysicalDeviceCopyMemoryIndirectFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceCopyMemoryIndirectFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    indirect_copy          Bool32
} 

// PhysicalDeviceCopyMemoryIndirectPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceCopyMemoryIndirectPropertiesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    supported_queues       QueueFlags
} 

type VkCmdCopyMemoryIndirectNV = fn (     C.CommandBuffer,     DeviceAddress,     u32,     u32) 

pub fn cmd_copy_memory_indirect_nv(
    command_buffer                                  C.CommandBuffer,
    copy_buffer_address                             DeviceAddress,
    copy_count                                      u32,
    stride                                          u32)  {
      f := VkCmdCopyMemoryIndirectNV((*loader_p).get_sym('vkCmdCopyMemoryIndirectNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyMemoryIndirectNV': ${err}")
        return 
    })
    f(
    command_buffer,
    copy_buffer_address,
    copy_count,
    stride)
}


type VkCmdCopyMemoryToImageIndirectNV = fn (     C.CommandBuffer,     DeviceAddress,     u32,     u32,     C.Image,     ImageLayout,     &ImageSubresourceLayers) 

pub fn cmd_copy_memory_to_image_indirect_nv(
    command_buffer                                  C.CommandBuffer,
    copy_buffer_address                             DeviceAddress,
    copy_count                                      u32,
    stride                                          u32,
    dst_image                                       C.Image,
    dst_image_layout                                ImageLayout,
    p_image_subresources                            &ImageSubresourceLayers)  {
      f := VkCmdCopyMemoryToImageIndirectNV((*loader_p).get_sym('vkCmdCopyMemoryToImageIndirectNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyMemoryToImageIndirectNV': ${err}")
        return 
    })
    f(
    command_buffer,
    copy_buffer_address,
    copy_count,
    stride,
    dst_image,
    dst_image_layout,
    p_image_subresources)
}




// VK_NV_memory_decompression is a preprocessor guard. Do not pass it to API calls.
const nv_memory_decompression = 1
pub const nv_memory_decompression_spec_version = 1
pub const nv_memory_decompression_extension_name = "VK_NV_memory_decompression"

// Flag bits for MemoryDecompressionMethodFlagBitsNV
pub type MemoryDecompressionMethodFlagBitsNV = u64
pub const memory_decompression_method_gdeflate_1_0_bit_nv = u64(0x00000001)


pub type MemoryDecompressionMethodFlagsNV = u64
pub struct DecompressMemoryRegionNV {
mut:
    src_address                               DeviceAddress
    dst_address                               DeviceAddress
    compressed_size                           DeviceSize
    decompressed_size                         DeviceSize
    decompression_method                      MemoryDecompressionMethodFlagsNV
} 

// PhysicalDeviceMemoryDecompressionFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMemoryDecompressionFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    memory_decompression   Bool32
} 

// PhysicalDeviceMemoryDecompressionPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceMemoryDecompressionPropertiesNV {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    decompression_methods                     MemoryDecompressionMethodFlagsNV
    max_decompression_indirect_count          u64
} 

type VkCmdDecompressMemoryNV = fn (     C.CommandBuffer,     u32,     &DecompressMemoryRegionNV) 

pub fn cmd_decompress_memory_nv(
    command_buffer                                  C.CommandBuffer,
    decompress_region_count                         u32,
    p_decompress_memory_regions                     &DecompressMemoryRegionNV)  {
      f := VkCmdDecompressMemoryNV((*loader_p).get_sym('vkCmdDecompressMemoryNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDecompressMemoryNV': ${err}")
        return 
    })
    f(
    command_buffer,
    decompress_region_count,
    p_decompress_memory_regions)
}


type VkCmdDecompressMemoryIndirectCountNV = fn (     C.CommandBuffer,     DeviceAddress,     DeviceAddress,     u32) 

pub fn cmd_decompress_memory_indirect_count_nv(
    command_buffer                                  C.CommandBuffer,
    indirect_commands_address                       DeviceAddress,
    indirect_commands_count_address                 DeviceAddress,
    stride                                          u32)  {
      f := VkCmdDecompressMemoryIndirectCountNV((*loader_p).get_sym('vkCmdDecompressMemoryIndirectCountNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDecompressMemoryIndirectCountNV': ${err}")
        return 
    })
    f(
    command_buffer,
    indirect_commands_address,
    indirect_commands_count_address,
    stride)
}




// VK_NV_device_generated_commands_compute is a preprocessor guard. Do not pass it to API calls.
const nv_device_generated_commands_compute = 1
pub const nv_device_generated_commands_compute_spec_version = 2
pub const nv_device_generated_commands_compute_extension_name = "VK_NV_device_generated_commands_compute"
// PhysicalDeviceDeviceGeneratedCommandsComputeFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDeviceGeneratedCommandsComputeFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_generated_compute Bool32
    device_generated_compute_pipelines Bool32
    device_generated_compute_capture_replay Bool32
} 

pub struct ComputePipelineIndirectBufferInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    device_address         DeviceAddress
    size                   DeviceSize
    pipeline_device_address_capture_replay DeviceAddress
} 

pub struct PipelineIndirectDeviceAddressInfoNV {
mut:
    s_type                     StructureType
    p_next                     voidptr
    pipeline_bind_point        PipelineBindPoint
    pipeline                   C.Pipeline
} 

pub struct BindPipelineIndirectCommandNV {
mut:
    pipeline_address       DeviceAddress
} 

type VkGetPipelineIndirectMemoryRequirementsNV = fn (     C.Device,     &ComputePipelineCreateInfo,     &MemoryRequirements2) 

pub fn get_pipeline_indirect_memory_requirements_nv(
    device                                          C.Device,
    p_create_info                                   &ComputePipelineCreateInfo,
    p_memory_requirements                           &MemoryRequirements2)  {
      f := VkGetPipelineIndirectMemoryRequirementsNV((*loader_p).get_sym('vkGetPipelineIndirectMemoryRequirementsNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetPipelineIndirectMemoryRequirementsNV': ${err}")
        return 
    })
    f(
    device,
    p_create_info,
    p_memory_requirements)
}


type VkCmdUpdatePipelineIndirectBufferNV = fn (     C.CommandBuffer,     PipelineBindPoint,     C.Pipeline) 

pub fn cmd_update_pipeline_indirect_buffer_nv(
    command_buffer                                  C.CommandBuffer,
    pipeline_bind_point                             PipelineBindPoint,
    pipeline                                        C.Pipeline)  {
      f := VkCmdUpdatePipelineIndirectBufferNV((*loader_p).get_sym('vkCmdUpdatePipelineIndirectBufferNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdUpdatePipelineIndirectBufferNV': ${err}")
        return 
    })
    f(
    command_buffer,
    pipeline_bind_point,
    pipeline)
}


type VkGetPipelineIndirectDeviceAddressNV = fn (     C.Device,     &PipelineIndirectDeviceAddressInfoNV) DeviceAddress

pub fn get_pipeline_indirect_device_address_nv(
    device                                          C.Device,
    p_info                                          &PipelineIndirectDeviceAddressInfoNV) DeviceAddress {
      f := VkGetPipelineIndirectDeviceAddressNV((*loader_p).get_sym("vkGetPipelineIndirectDeviceAddressNV"
    ) or { 
        panic("Couldn't load symbol for 'vkGetPipelineIndirectDeviceAddressNV': ${err}") })
    return f(
    device,
    p_info)
}




// VK_NV_linear_color_attachment is a preprocessor guard. Do not pass it to API calls.
const nv_linear_color_attachment = 1
pub const nv_linear_color_attachment_spec_version = 1
pub const nv_linear_color_attachment_extension_name = "VK_NV_linear_color_attachment"
// PhysicalDeviceLinearColorAttachmentFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceLinearColorAttachmentFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    linear_color_attachment Bool32
} 



// VK_GOOGLE_surfaceless_query is a preprocessor guard. Do not pass it to API calls.
const google_surfaceless_query = 1
pub const google_surfaceless_query_spec_version = 2
pub const google_surfaceless_query_extension_name = "VK_GOOGE_surfaceless_query"


// VK_EXT_image_compression_control_swapchain is a preprocessor guard. Do not pass it to API calls.
const ext_image_compression_control_swapchain = 1
pub const ext_image_compression_control_swapchain_spec_version = 1
pub const ext_image_compression_control_swapchain_extension_name = "VK_EXT_image_compression_control_swapchain"
// PhysicalDeviceImageCompressionControlSwapchainFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceImageCompressionControlSwapchainFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    image_compression_control_swapchain Bool32
} 



// VK_QCOM_image_processing is a preprocessor guard. Do not pass it to API calls.
const qcom_image_processing = 1
pub const qcom_image_processing_spec_version = 1
pub const qcom_image_processing_extension_name = "VK_QCOM_image_processing"
// ImageViewSampleWeightCreateInfoQCOM extends VkImageViewCreateInfo
pub struct ImageViewSampleWeightCreateInfoQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    filter_center          Offset2D
    filter_size            Extent2D
    num_phases             u32
} 

// PhysicalDeviceImageProcessingFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceImageProcessingFeaturesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    texture_sample_weighted Bool32
    texture_box_filter     Bool32
    texture_block_match    Bool32
} 

// PhysicalDeviceImageProcessingPropertiesQCOM extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceImageProcessingPropertiesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_weight_filter_phases u32
    max_weight_filter_dimension Extent2D
    max_block_match_region Extent2D
    max_box_filter_block_size Extent2D
} 



// VK_EXT_nested_command_buffer is a preprocessor guard. Do not pass it to API calls.
const ext_nested_command_buffer = 1
pub const ext_nested_command_buffer_spec_version = 1
pub const ext_nested_command_buffer_extension_name = "VK_EXT_nested_command_buffer"
// PhysicalDeviceNestedCommandBufferFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceNestedCommandBufferFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    nested_command_buffer  Bool32
    nested_command_buffer_rendering Bool32
    nested_command_buffer_simultaneous_use Bool32
} 

// PhysicalDeviceNestedCommandBufferPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceNestedCommandBufferPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_command_buffer_nesting_level u32
} 



// VK_EXT_external_memory_acquire_unmodified is a preprocessor guard. Do not pass it to API calls.
const ext_external_memory_acquire_unmodified = 1
pub const ext_external_memory_acquire_unmodified_spec_version = 1
pub const ext_external_memory_acquire_unmodified_extension_name = "VK_EXT_external_memory_acquire_unmodified"
// ExternalMemoryAcquireUnmodifiedEXT extends VkBufferMemoryBarrier,VkBufferMemoryBarrier2,VkImageMemoryBarrier,VkImageMemoryBarrier2
pub struct ExternalMemoryAcquireUnmodifiedEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    acquire_unmodified_memory Bool32
} 



// VK_EXT_extended_dynamic_state3 is a preprocessor guard. Do not pass it to API calls.
const ext_extended_dynamic_state3 = 1
pub const ext_extended_dynamic_state_3_spec_version = 2
pub const ext_extended_dynamic_state_3_extension_name = "VK_EXT_extended_dynamic_state3"
// PhysicalDeviceExtendedDynamicState3FeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceExtendedDynamicState3FeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    extended_dynamic_state3_tessellation_domain_origin Bool32
    extended_dynamic_state3_depth_clamp_enable Bool32
    extended_dynamic_state3_polygon_mode Bool32
    extended_dynamic_state3_rasterization_samples Bool32
    extended_dynamic_state3_sample_mask Bool32
    extended_dynamic_state3_alpha_to_coverage_enable Bool32
    extended_dynamic_state3_alpha_to_one_enable Bool32
    extended_dynamic_state3_logic_op_enable Bool32
    extended_dynamic_state3_color_blend_enable Bool32
    extended_dynamic_state3_color_blend_equation Bool32
    extended_dynamic_state3_color_write_mask Bool32
    extended_dynamic_state3_rasterization_stream Bool32
    extended_dynamic_state3_conservative_rasterization_mode Bool32
    extended_dynamic_state3_extra_primitive_overestimation_size Bool32
    extended_dynamic_state3_depth_clip_enable Bool32
    extended_dynamic_state3_sample_locations_enable Bool32
    extended_dynamic_state3_color_blend_advanced Bool32
    extended_dynamic_state3_provoking_vertex_mode Bool32
    extended_dynamic_state3_line_rasterization_mode Bool32
    extended_dynamic_state3_line_stipple_enable Bool32
    extended_dynamic_state3_depth_clip_negative_one_to_one Bool32
    extended_dynamic_state3_viewport_w_scaling_enable Bool32
    extended_dynamic_state3_viewport_swizzle Bool32
    extended_dynamic_state3_coverage_to_color_enable Bool32
    extended_dynamic_state3_coverage_to_color_location Bool32
    extended_dynamic_state3_coverage_modulation_mode Bool32
    extended_dynamic_state3_coverage_modulation_table_enable Bool32
    extended_dynamic_state3_coverage_modulation_table Bool32
    extended_dynamic_state3_coverage_reduction_mode Bool32
    extended_dynamic_state3_representative_fragment_test_enable Bool32
    extended_dynamic_state3_shading_rate_image_enable Bool32
} 

// PhysicalDeviceExtendedDynamicState3PropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceExtendedDynamicState3PropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    dynamic_primitive_topology_unrestricted Bool32
} 

pub struct ColorBlendEquationEXT {
mut:
    src_color_blend_factor BlendFactor
    dst_color_blend_factor BlendFactor
    color_blend_op       BlendOp
    src_alpha_blend_factor BlendFactor
    dst_alpha_blend_factor BlendFactor
    alpha_blend_op       BlendOp
} 

pub struct ColorBlendAdvancedEXT {
mut:
    advanced_blend_op        BlendOp
    src_premultiplied        Bool32
    dst_premultiplied        Bool32
    blend_overlap            BlendOverlapEXT
    clamp_results            Bool32
} 

type VkCmdSetTessellationDomainOriginEXT = fn (     C.CommandBuffer,     TessellationDomainOrigin) 

pub fn cmd_set_tessellation_domain_origin_ext(
    command_buffer                                  C.CommandBuffer,
    domain_origin                                   TessellationDomainOrigin)  {
      f := VkCmdSetTessellationDomainOriginEXT((*loader_p).get_sym('vkCmdSetTessellationDomainOriginEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetTessellationDomainOriginEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    domain_origin)
}


type VkCmdSetDepthClampEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_depth_clamp_enable_ext(
    command_buffer                                  C.CommandBuffer,
    depth_clamp_enable                              Bool32)  {
      f := VkCmdSetDepthClampEnableEXT((*loader_p).get_sym('vkCmdSetDepthClampEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthClampEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_clamp_enable)
}


type VkCmdSetPolygonModeEXT = fn (     C.CommandBuffer,     PolygonMode) 

pub fn cmd_set_polygon_mode_ext(
    command_buffer                                  C.CommandBuffer,
    polygon_mode                                    PolygonMode)  {
      f := VkCmdSetPolygonModeEXT((*loader_p).get_sym('vkCmdSetPolygonModeEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetPolygonModeEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    polygon_mode)
}


type VkCmdSetRasterizationSamplesEXT = fn (     C.CommandBuffer,     SampleCountFlagBits) 

pub fn cmd_set_rasterization_samples_ext(
    command_buffer                                  C.CommandBuffer,
    rasterization_samples                           SampleCountFlagBits)  {
      f := VkCmdSetRasterizationSamplesEXT((*loader_p).get_sym('vkCmdSetRasterizationSamplesEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetRasterizationSamplesEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    rasterization_samples)
}


type VkCmdSetSampleMaskEXT = fn (     C.CommandBuffer,     SampleCountFlagBits,     &SampleMask) 

pub fn cmd_set_sample_mask_ext(
    command_buffer                                  C.CommandBuffer,
    samples                                         SampleCountFlagBits,
    p_sample_mask                                   &SampleMask)  {
      f := VkCmdSetSampleMaskEXT((*loader_p).get_sym('vkCmdSetSampleMaskEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetSampleMaskEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    samples,
    p_sample_mask)
}


type VkCmdSetAlphaToCoverageEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_alpha_to_coverage_enable_ext(
    command_buffer                                  C.CommandBuffer,
    alpha_to_coverage_enable                        Bool32)  {
      f := VkCmdSetAlphaToCoverageEnableEXT((*loader_p).get_sym('vkCmdSetAlphaToCoverageEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetAlphaToCoverageEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    alpha_to_coverage_enable)
}


type VkCmdSetAlphaToOneEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_alpha_to_one_enable_ext(
    command_buffer                                  C.CommandBuffer,
    alpha_to_one_enable                             Bool32)  {
      f := VkCmdSetAlphaToOneEnableEXT((*loader_p).get_sym('vkCmdSetAlphaToOneEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetAlphaToOneEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    alpha_to_one_enable)
}


type VkCmdSetLogicOpEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_logic_op_enable_ext(
    command_buffer                                  C.CommandBuffer,
    logic_op_enable                                 Bool32)  {
      f := VkCmdSetLogicOpEnableEXT((*loader_p).get_sym('vkCmdSetLogicOpEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetLogicOpEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    logic_op_enable)
}


type VkCmdSetColorBlendEnableEXT = fn (     C.CommandBuffer,     u32,     u32,     &Bool32) 

pub fn cmd_set_color_blend_enable_ext(
    command_buffer                                  C.CommandBuffer,
    first_attachment                                u32,
    attachment_count                                u32,
    p_color_blend_enables                           &Bool32)  {
      f := VkCmdSetColorBlendEnableEXT((*loader_p).get_sym('vkCmdSetColorBlendEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetColorBlendEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    first_attachment,
    attachment_count,
    p_color_blend_enables)
}


type VkCmdSetColorBlendEquationEXT = fn (     C.CommandBuffer,     u32,     u32,     &ColorBlendEquationEXT) 

pub fn cmd_set_color_blend_equation_ext(
    command_buffer                                  C.CommandBuffer,
    first_attachment                                u32,
    attachment_count                                u32,
    p_color_blend_equations                         &ColorBlendEquationEXT)  {
      f := VkCmdSetColorBlendEquationEXT((*loader_p).get_sym('vkCmdSetColorBlendEquationEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetColorBlendEquationEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    first_attachment,
    attachment_count,
    p_color_blend_equations)
}


type VkCmdSetColorWriteMaskEXT = fn (     C.CommandBuffer,     u32,     u32,     &ColorComponentFlags) 

pub fn cmd_set_color_write_mask_ext(
    command_buffer                                  C.CommandBuffer,
    first_attachment                                u32,
    attachment_count                                u32,
    p_color_write_masks                             &ColorComponentFlags)  {
      f := VkCmdSetColorWriteMaskEXT((*loader_p).get_sym('vkCmdSetColorWriteMaskEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetColorWriteMaskEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    first_attachment,
    attachment_count,
    p_color_write_masks)
}


type VkCmdSetRasterizationStreamEXT = fn (     C.CommandBuffer,     u32) 

pub fn cmd_set_rasterization_stream_ext(
    command_buffer                                  C.CommandBuffer,
    rasterization_stream                            u32)  {
      f := VkCmdSetRasterizationStreamEXT((*loader_p).get_sym('vkCmdSetRasterizationStreamEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetRasterizationStreamEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    rasterization_stream)
}


type VkCmdSetConservativeRasterizationModeEXT = fn (     C.CommandBuffer,     ConservativeRasterizationModeEXT) 

pub fn cmd_set_conservative_rasterization_mode_ext(
    command_buffer                                  C.CommandBuffer,
    conservative_rasterization_mode                 ConservativeRasterizationModeEXT)  {
      f := VkCmdSetConservativeRasterizationModeEXT((*loader_p).get_sym('vkCmdSetConservativeRasterizationModeEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetConservativeRasterizationModeEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    conservative_rasterization_mode)
}


type VkCmdSetExtraPrimitiveOverestimationSizeEXT = fn (     C.CommandBuffer,     f32) 

pub fn cmd_set_extra_primitive_overestimation_size_ext(
    command_buffer                                  C.CommandBuffer,
    extra_primitive_overestimation_size             f32)  {
      f := VkCmdSetExtraPrimitiveOverestimationSizeEXT((*loader_p).get_sym('vkCmdSetExtraPrimitiveOverestimationSizeEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetExtraPrimitiveOverestimationSizeEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    extra_primitive_overestimation_size)
}


type VkCmdSetDepthClipEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_depth_clip_enable_ext(
    command_buffer                                  C.CommandBuffer,
    depth_clip_enable                               Bool32)  {
      f := VkCmdSetDepthClipEnableEXT((*loader_p).get_sym('vkCmdSetDepthClipEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthClipEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    depth_clip_enable)
}


type VkCmdSetSampleLocationsEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_sample_locations_enable_ext(
    command_buffer                                  C.CommandBuffer,
    sample_locations_enable                         Bool32)  {
      f := VkCmdSetSampleLocationsEnableEXT((*loader_p).get_sym('vkCmdSetSampleLocationsEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetSampleLocationsEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    sample_locations_enable)
}


type VkCmdSetColorBlendAdvancedEXT = fn (     C.CommandBuffer,     u32,     u32,     &ColorBlendAdvancedEXT) 

pub fn cmd_set_color_blend_advanced_ext(
    command_buffer                                  C.CommandBuffer,
    first_attachment                                u32,
    attachment_count                                u32,
    p_color_blend_advanced                          &ColorBlendAdvancedEXT)  {
      f := VkCmdSetColorBlendAdvancedEXT((*loader_p).get_sym('vkCmdSetColorBlendAdvancedEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetColorBlendAdvancedEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    first_attachment,
    attachment_count,
    p_color_blend_advanced)
}


type VkCmdSetProvokingVertexModeEXT = fn (     C.CommandBuffer,     ProvokingVertexModeEXT) 

pub fn cmd_set_provoking_vertex_mode_ext(
    command_buffer                                  C.CommandBuffer,
    provoking_vertex_mode                           ProvokingVertexModeEXT)  {
      f := VkCmdSetProvokingVertexModeEXT((*loader_p).get_sym('vkCmdSetProvokingVertexModeEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetProvokingVertexModeEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    provoking_vertex_mode)
}


type VkCmdSetLineRasterizationModeEXT = fn (     C.CommandBuffer,     LineRasterizationModeEXT) 

pub fn cmd_set_line_rasterization_mode_ext(
    command_buffer                                  C.CommandBuffer,
    line_rasterization_mode                         LineRasterizationModeEXT)  {
      f := VkCmdSetLineRasterizationModeEXT((*loader_p).get_sym('vkCmdSetLineRasterizationModeEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetLineRasterizationModeEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    line_rasterization_mode)
}


type VkCmdSetLineStippleEnableEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_line_stipple_enable_ext(
    command_buffer                                  C.CommandBuffer,
    stippled_line_enable                            Bool32)  {
      f := VkCmdSetLineStippleEnableEXT((*loader_p).get_sym('vkCmdSetLineStippleEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetLineStippleEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    stippled_line_enable)
}


type VkCmdSetDepthClipNegativeOneToOneEXT = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_depth_clip_negative_one_to_one_ext(
    command_buffer                                  C.CommandBuffer,
    negative_one_to_one                             Bool32)  {
      f := VkCmdSetDepthClipNegativeOneToOneEXT((*loader_p).get_sym('vkCmdSetDepthClipNegativeOneToOneEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetDepthClipNegativeOneToOneEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    negative_one_to_one)
}


type VkCmdSetViewportWScalingEnableNV = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_viewport_w_scaling_enable_nv(
    command_buffer                                  C.CommandBuffer,
    viewport_w_scaling_enable                       Bool32)  {
      f := VkCmdSetViewportWScalingEnableNV((*loader_p).get_sym('vkCmdSetViewportWScalingEnableNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetViewportWScalingEnableNV': ${err}")
        return 
    })
    f(
    command_buffer,
    viewport_w_scaling_enable)
}


type VkCmdSetViewportSwizzleNV = fn (     C.CommandBuffer,     u32,     u32,     &ViewportSwizzleNV) 

pub fn cmd_set_viewport_swizzle_nv(
    command_buffer                                  C.CommandBuffer,
    first_viewport                                  u32,
    viewport_count                                  u32,
    p_viewport_swizzles                             &ViewportSwizzleNV)  {
      f := VkCmdSetViewportSwizzleNV((*loader_p).get_sym('vkCmdSetViewportSwizzleNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetViewportSwizzleNV': ${err}")
        return 
    })
    f(
    command_buffer,
    first_viewport,
    viewport_count,
    p_viewport_swizzles)
}


type VkCmdSetCoverageToColorEnableNV = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_coverage_to_color_enable_nv(
    command_buffer                                  C.CommandBuffer,
    coverage_to_color_enable                        Bool32)  {
      f := VkCmdSetCoverageToColorEnableNV((*loader_p).get_sym('vkCmdSetCoverageToColorEnableNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetCoverageToColorEnableNV': ${err}")
        return 
    })
    f(
    command_buffer,
    coverage_to_color_enable)
}


type VkCmdSetCoverageToColorLocationNV = fn (     C.CommandBuffer,     u32) 

pub fn cmd_set_coverage_to_color_location_nv(
    command_buffer                                  C.CommandBuffer,
    coverage_to_color_location                      u32)  {
      f := VkCmdSetCoverageToColorLocationNV((*loader_p).get_sym('vkCmdSetCoverageToColorLocationNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetCoverageToColorLocationNV': ${err}")
        return 
    })
    f(
    command_buffer,
    coverage_to_color_location)
}


type VkCmdSetCoverageModulationModeNV = fn (     C.CommandBuffer,     CoverageModulationModeNV) 

pub fn cmd_set_coverage_modulation_mode_nv(
    command_buffer                                  C.CommandBuffer,
    coverage_modulation_mode                        CoverageModulationModeNV)  {
      f := VkCmdSetCoverageModulationModeNV((*loader_p).get_sym('vkCmdSetCoverageModulationModeNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetCoverageModulationModeNV': ${err}")
        return 
    })
    f(
    command_buffer,
    coverage_modulation_mode)
}


type VkCmdSetCoverageModulationTableEnableNV = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_coverage_modulation_table_enable_nv(
    command_buffer                                  C.CommandBuffer,
    coverage_modulation_table_enable                Bool32)  {
      f := VkCmdSetCoverageModulationTableEnableNV((*loader_p).get_sym('vkCmdSetCoverageModulationTableEnableNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetCoverageModulationTableEnableNV': ${err}")
        return 
    })
    f(
    command_buffer,
    coverage_modulation_table_enable)
}


type VkCmdSetCoverageModulationTableNV = fn (     C.CommandBuffer,     u32,     &f32) 

pub fn cmd_set_coverage_modulation_table_nv(
    command_buffer                                  C.CommandBuffer,
    coverage_modulation_table_count                 u32,
    p_coverage_modulation_table                     &f32)  {
      f := VkCmdSetCoverageModulationTableNV((*loader_p).get_sym('vkCmdSetCoverageModulationTableNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetCoverageModulationTableNV': ${err}")
        return 
    })
    f(
    command_buffer,
    coverage_modulation_table_count,
    p_coverage_modulation_table)
}


type VkCmdSetShadingRateImageEnableNV = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_shading_rate_image_enable_nv(
    command_buffer                                  C.CommandBuffer,
    shading_rate_image_enable                       Bool32)  {
      f := VkCmdSetShadingRateImageEnableNV((*loader_p).get_sym('vkCmdSetShadingRateImageEnableNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetShadingRateImageEnableNV': ${err}")
        return 
    })
    f(
    command_buffer,
    shading_rate_image_enable)
}


type VkCmdSetRepresentativeFragmentTestEnableNV = fn (     C.CommandBuffer,     Bool32) 

pub fn cmd_set_representative_fragment_test_enable_nv(
    command_buffer                                  C.CommandBuffer,
    representative_fragment_test_enable             Bool32)  {
      f := VkCmdSetRepresentativeFragmentTestEnableNV((*loader_p).get_sym('vkCmdSetRepresentativeFragmentTestEnableNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetRepresentativeFragmentTestEnableNV': ${err}")
        return 
    })
    f(
    command_buffer,
    representative_fragment_test_enable)
}


type VkCmdSetCoverageReductionModeNV = fn (     C.CommandBuffer,     CoverageReductionModeNV) 

pub fn cmd_set_coverage_reduction_mode_nv(
    command_buffer                                  C.CommandBuffer,
    coverage_reduction_mode                         CoverageReductionModeNV)  {
      f := VkCmdSetCoverageReductionModeNV((*loader_p).get_sym('vkCmdSetCoverageReductionModeNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetCoverageReductionModeNV': ${err}")
        return 
    })
    f(
    command_buffer,
    coverage_reduction_mode)
}




// VK_EXT_subpass_merge_feedback is a preprocessor guard. Do not pass it to API calls.
const ext_subpass_merge_feedback = 1
pub const ext_subpass_merge_feedback_spec_version = 2
pub const ext_subpass_merge_feedback_extension_name = "VK_EXT_subpass_merge_feedback"

pub enum SubpassMergeStatusEXT {
    subpass_merge_status_merged_ext = int(0)
    subpass_merge_status_disallowed_ext = int(1)
    subpass_merge_status_not_merged_side_effects_ext = int(2)
    subpass_merge_status_not_merged_samples_mismatch_ext = int(3)
    subpass_merge_status_not_merged_views_mismatch_ext = int(4)
    subpass_merge_status_not_merged_aliasing_ext = int(5)
    subpass_merge_status_not_merged_dependencies_ext = int(6)
    subpass_merge_status_not_merged_incompatible_input_attachment_ext = int(7)
    subpass_merge_status_not_merged_too_many_attachments_ext = int(8)
    subpass_merge_status_not_merged_insufficient_storage_ext = int(9)
    subpass_merge_status_not_merged_depth_stencil_count_ext = int(10)
    subpass_merge_status_not_merged_resolve_attachment_reuse_ext = int(11)
    subpass_merge_status_not_merged_single_subpass_ext = int(12)
    subpass_merge_status_not_merged_unspecified_ext = int(13)
    subpass_merge_status_max_enum_ext = int(0x7FFFFFFF)
}

// PhysicalDeviceSubpassMergeFeedbackFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceSubpassMergeFeedbackFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    subpass_merge_feedback Bool32
} 

// RenderPassCreationControlEXT extends VkRenderPassCreateInfo2,VkSubpassDescription2
pub struct RenderPassCreationControlEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    disallow_merging       Bool32
} 

pub struct RenderPassCreationFeedbackInfoEXT {
mut:
    post_merge_subpass_count u32
} 

// RenderPassCreationFeedbackCreateInfoEXT extends VkRenderPassCreateInfo2
pub struct RenderPassCreationFeedbackCreateInfoEXT {
mut:
    s_type                                      StructureType
    p_next                                      voidptr
    p_render_pass_feedback                      &RenderPassCreationFeedbackInfoEXT
} 

pub struct RenderPassSubpassFeedbackInfoEXT {
mut:
    subpass_merge_status           SubpassMergeStatusEXT
    description                    []char
    post_merge_index               u32
} 

// RenderPassSubpassFeedbackCreateInfoEXT extends VkSubpassDescription2
pub struct RenderPassSubpassFeedbackCreateInfoEXT {
mut:
    s_type                                     StructureType
    p_next                                     voidptr
    p_subpass_feedback                         &RenderPassSubpassFeedbackInfoEXT
} 



// VK_LUNARG_direct_driver_loading is a preprocessor guard. Do not pass it to API calls.
const lunarg_direct_driver_loading = 1
pub const lunarg_direct_driver_loading_spec_version = 1
pub const lunarg_direct_driver_loading_extension_name = "VK_NARG_direct_driver_loading"

pub enum DirectDriverLoadingModeLUNARG {
    direct_driver_loading_mode_exclusive_lunarg = int(0)
    direct_driver_loading_mode_inclusive_lunarg = int(1)
    direct_driver_loading_mode_max_enum_lunarg = int(0x7FFFFFFF)
}

pub type DirectDriverLoadingFlagsLUNARG = u32
pub type PFN_vkGetInstanceProcAddrLUNARG = fn (   instanceconst                     C.Instance,   pName                             &char) voidptr
pub struct DirectDriverLoadingInfoLUNARG {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    flags                                   DirectDriverLoadingFlagsLUNARG
    pfn_get_instance_proc_addr              PFN_vkGetInstanceProcAddrLUNARG = unsafe { nil }
} 

// DirectDriverLoadingListLUNARG extends VkInstanceCreateInfo
pub struct DirectDriverLoadingListLUNARG {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    mode                                          DirectDriverLoadingModeLUNARG
    driver_count                                  u32
    p_drivers                                     &DirectDriverLoadingInfoLUNARG
} 



// VK_EXT_shader_module_identifier is a preprocessor guard. Do not pass it to API calls.
const ext_shader_module_identifier = 1
pub const max_shader_module_identifier_size_ext = u32(32)
pub const ext_shader_module_identifier_spec_version = 1
pub const ext_shader_module_identifier_extension_name = "VK_EXT_shader_module_identifier"
// PhysicalDeviceShaderModuleIdentifierFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderModuleIdentifierFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_module_identifier Bool32
} 

// PhysicalDeviceShaderModuleIdentifierPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceShaderModuleIdentifierPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_module_identifier_algorithm_uuid []u8
} 

// PipelineShaderStageModuleIdentifierCreateInfoEXT extends VkPipelineShaderStageCreateInfo
pub struct PipelineShaderStageModuleIdentifierCreateInfoEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    identifier_size        u32
    p_identifier           &u8
} 

pub struct ShaderModuleIdentifierEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    identifier_size        u32
    identifier             []u8
} 

type VkGetShaderModuleIdentifierEXT = fn (     C.Device,     C.ShaderModule,     &ShaderModuleIdentifierEXT) 

pub fn get_shader_module_identifier_ext(
    device                                          C.Device,
    shader_module                                   C.ShaderModule,
    p_identifier                                    &ShaderModuleIdentifierEXT)  {
      f := VkGetShaderModuleIdentifierEXT((*loader_p).get_sym('vkGetShaderModuleIdentifierEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetShaderModuleIdentifierEXT': ${err}")
        return 
    })
    f(
    device,
    shader_module,
    p_identifier)
}


type VkGetShaderModuleCreateInfoIdentifierEXT = fn (     C.Device,     &ShaderModuleCreateInfo,     &ShaderModuleIdentifierEXT) 

pub fn get_shader_module_create_info_identifier_ext(
    device                                          C.Device,
    p_create_info                                   &ShaderModuleCreateInfo,
    p_identifier                                    &ShaderModuleIdentifierEXT)  {
      f := VkGetShaderModuleCreateInfoIdentifierEXT((*loader_p).get_sym('vkGetShaderModuleCreateInfoIdentifierEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetShaderModuleCreateInfoIdentifierEXT': ${err}")
        return 
    })
    f(
    device,
    p_create_info,
    p_identifier)
}




// VK_EXT_rasterization_order_attachment_access is a preprocessor guard. Do not pass it to API calls.
const ext_rasterization_order_attachment_access = 1
pub const ext_rasterization_order_attachment_access_spec_version = 1
pub const ext_rasterization_order_attachment_access_extension_name = "VK_EXT_rasterization_order_attachment_access"


// VK_NV_optical_flow is a preprocessor guard. Do not pass it to API calls.
const nv_optical_flow = 1
pub type C.OpticalFlowSessionNV = voidptr
pub const nv_optical_flow_spec_version      = 1
pub const nv_optical_flow_extension_name    = "VK_NV_optical_flow"

pub enum OpticalFlowPerformanceLevelNV {
    optical_flow_performance_level_unknown_nv = int(0)
    optical_flow_performance_level_slow_nv = int(1)
    optical_flow_performance_level_medium_nv = int(2)
    optical_flow_performance_level_fast_nv = int(3)
    optical_flow_performance_level_max_enum_nv = int(0x7FFFFFFF)
}


pub enum OpticalFlowSessionBindingPointNV {
    optical_flow_session_binding_point_unknown_nv = int(0)
    optical_flow_session_binding_point_input_nv = int(1)
    optical_flow_session_binding_point_reference_nv = int(2)
    optical_flow_session_binding_point_hint_nv = int(3)
    optical_flow_session_binding_point_flow_vector_nv = int(4)
    optical_flow_session_binding_point_backward_flow_vector_nv = int(5)
    optical_flow_session_binding_point_cost_nv = int(6)
    optical_flow_session_binding_point_backward_cost_nv = int(7)
    optical_flow_session_binding_point_global_flow_nv = int(8)
    optical_flow_session_binding_point_max_enum_nv = int(0x7FFFFFFF)
}


pub enum OpticalFlowGridSizeFlagBitsNV {
    optical_flow_grid_size_unknown_nv = int(0)
    optical_flow_grid_size_1x1_bit_nv = int(0x00000001)
    optical_flow_grid_size_2x2_bit_nv = int(0x00000002)
    optical_flow_grid_size_4x4_bit_nv = int(0x00000004)
    optical_flow_grid_size_8x8_bit_nv = int(0x00000008)
    optical_flow_grid_size_flag_bits_max_enum_nv = int(0x7FFFFFFF)
}

pub type OpticalFlowGridSizeFlagsNV = u32

pub enum OpticalFlowUsageFlagBitsNV {
    optical_flow_usage_unknown_nv = int(0)
    optical_flow_usage_input_bit_nv = int(0x00000001)
    optical_flow_usage_output_bit_nv = int(0x00000002)
    optical_flow_usage_hint_bit_nv = int(0x00000004)
    optical_flow_usage_cost_bit_nv = int(0x00000008)
    optical_flow_usage_global_flow_bit_nv = int(0x00000010)
    optical_flow_usage_flag_bits_max_enum_nv = int(0x7FFFFFFF)
}

pub type OpticalFlowUsageFlagsNV = u32

pub enum OpticalFlowSessionCreateFlagBitsNV {
    optical_flow_session_create_enable_hint_bit_nv = int(0x00000001)
    optical_flow_session_create_enable_cost_bit_nv = int(0x00000002)
    optical_flow_session_create_enable_global_flow_bit_nv = int(0x00000004)
    optical_flow_session_create_allow_regions_bit_nv = int(0x00000008)
    optical_flow_session_create_both_directions_bit_nv = int(0x00000010)
    optical_flow_session_create_flag_bits_max_enum_nv = int(0x7FFFFFFF)
}

pub type OpticalFlowSessionCreateFlagsNV = u32

pub enum OpticalFlowExecuteFlagBitsNV {
    optical_flow_execute_disable_temporal_hints_bit_nv = int(0x00000001)
    optical_flow_execute_flag_bits_max_enum_nv = int(0x7FFFFFFF)
}

pub type OpticalFlowExecuteFlagsNV = u32
// PhysicalDeviceOpticalFlowFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceOpticalFlowFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    optical_flow           Bool32
} 

// PhysicalDeviceOpticalFlowPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceOpticalFlowPropertiesNV {
mut:
    s_type                              StructureType
    p_next                              voidptr
    supported_output_grid_sizes         OpticalFlowGridSizeFlagsNV
    supported_hint_grid_sizes           OpticalFlowGridSizeFlagsNV
    hint_supported                      Bool32
    cost_supported                      Bool32
    bidirectional_flow_supported        Bool32
    global_flow_supported               Bool32
    min_width                           u32
    min_height                          u32
    max_width                           u32
    max_height                          u32
    max_num_regions_of_interest         u32
} 

// OpticalFlowImageFormatInfoNV extends VkPhysicalDeviceImageFormatInfo2,VkImageCreateInfo
pub struct OpticalFlowImageFormatInfoNV {
mut:
    s_type                           StructureType
    p_next                           voidptr
    usage                            OpticalFlowUsageFlagsNV
} 

pub struct OpticalFlowImageFormatPropertiesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    format                 Format
} 

pub struct OpticalFlowSessionCreateInfoNV {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    width                                    u32
    height                                   u32
    image_format                             Format
    flow_vector_format                       Format
    cost_format                              Format
    output_grid_size                         OpticalFlowGridSizeFlagsNV
    hint_grid_size                           OpticalFlowGridSizeFlagsNV
    performance_level                        OpticalFlowPerformanceLevelNV
    flags                                    OpticalFlowSessionCreateFlagsNV
} 

// OpticalFlowSessionCreatePrivateDataInfoNV extends VkOpticalFlowSessionCreateInfoNV
pub struct OpticalFlowSessionCreatePrivateDataInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    id                     u32
    size                   u32
    p_private_data         voidptr
} 

pub struct OpticalFlowExecuteInfoNV {
mut:
    s_type                             StructureType
    p_next                             voidptr
    flags                              OpticalFlowExecuteFlagsNV
    region_count                       u32
    p_regions                          &Rect2D
} 

type VkGetPhysicalDeviceOpticalFlowImageFormatsNV = fn (     C.PhysicalDevice,     &OpticalFlowImageFormatInfoNV,     &u32,     &OpticalFlowImageFormatPropertiesNV) Result

pub fn get_physical_device_optical_flow_image_formats_nv(
    physical_device                                 C.PhysicalDevice,
    p_optical_flow_image_format_info                &OpticalFlowImageFormatInfoNV,
    p_format_count                                  &u32,
    p_image_format_properties                       &OpticalFlowImageFormatPropertiesNV) Result {
      f := VkGetPhysicalDeviceOpticalFlowImageFormatsNV((*loader_p).get_sym('vkGetPhysicalDeviceOpticalFlowImageFormatsNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetPhysicalDeviceOpticalFlowImageFormatsNV': ${err}")
        return Result.error_unknown
    })
    return f(
    physical_device,
    p_optical_flow_image_format_info,
    p_format_count,
    p_image_format_properties)
}


type VkCreateOpticalFlowSessionNV = fn (     C.Device,     &OpticalFlowSessionCreateInfoNV,     &AllocationCallbacks,     &C.OpticalFlowSessionNV) Result

pub fn create_optical_flow_session_nv(
    device                                          C.Device,
    p_create_info                                   &OpticalFlowSessionCreateInfoNV,
    p_allocator                                     &AllocationCallbacks,
    p_session                                       &C.OpticalFlowSessionNV) Result {
      f := VkCreateOpticalFlowSessionNV((*loader_p).get_sym('vkCreateOpticalFlowSessionNV'
    ) or { 
        println("Couldn't load symbol for 'vkCreateOpticalFlowSessionNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_session)
}


type VkDestroyOpticalFlowSessionNV = fn (     C.Device,     C.OpticalFlowSessionNV,     &AllocationCallbacks) 

pub fn destroy_optical_flow_session_nv(
    device                                          C.Device,
    session                                         C.OpticalFlowSessionNV,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyOpticalFlowSessionNV((*loader_p).get_sym('vkDestroyOpticalFlowSessionNV'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyOpticalFlowSessionNV': ${err}")
        return 
    })
    f(
    device,
    session,
    p_allocator)
}


type VkBindOpticalFlowSessionImageNV = fn (     C.Device,     C.OpticalFlowSessionNV,     OpticalFlowSessionBindingPointNV,     C.ImageView,     ImageLayout) Result

pub fn bind_optical_flow_session_image_nv(
    device                                          C.Device,
    session                                         C.OpticalFlowSessionNV,
    binding_point                                   OpticalFlowSessionBindingPointNV,
    view                                            C.ImageView,
    layout                                          ImageLayout) Result {
      f := VkBindOpticalFlowSessionImageNV((*loader_p).get_sym('vkBindOpticalFlowSessionImageNV'
    ) or { 
        println("Couldn't load symbol for 'vkBindOpticalFlowSessionImageNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    session,
    binding_point,
    view,
    layout)
}


type VkCmdOpticalFlowExecuteNV = fn (     C.CommandBuffer,     C.OpticalFlowSessionNV,     &OpticalFlowExecuteInfoNV) 

pub fn cmd_optical_flow_execute_nv(
    command_buffer                                  C.CommandBuffer,
    session                                         C.OpticalFlowSessionNV,
    p_execute_info                                  &OpticalFlowExecuteInfoNV)  {
      f := VkCmdOpticalFlowExecuteNV((*loader_p).get_sym('vkCmdOpticalFlowExecuteNV'
    ) or { 
        println("Couldn't load symbol for 'vkCmdOpticalFlowExecuteNV': ${err}")
        return 
    })
    f(
    command_buffer,
    session,
    p_execute_info)
}




// VK_EXT_legacy_dithering is a preprocessor guard. Do not pass it to API calls.
const ext_legacy_dithering = 1
pub const ext_legacy_dithering_spec_version = 1
pub const ext_legacy_dithering_extension_name = "VK_EXT_legacy_dithering"
// PhysicalDeviceLegacyDitheringFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceLegacyDitheringFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    legacy_dithering       Bool32
} 



// VK_EXT_pipeline_protected_access is a preprocessor guard. Do not pass it to API calls.
const ext_pipeline_protected_access = 1
pub const ext_pipeline_protected_access_spec_version = 1
pub const ext_pipeline_protected_access_extension_name = "VK_EXT_pipeline_protected_access"
// PhysicalDevicePipelineProtectedAccessFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePipelineProtectedAccessFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pipeline_protected_access Bool32
} 



// VK_ANDROID_external_format_resolve is a preprocessor guard. Do not pass it to API calls.
const android_external_format_resolve = 1
pub const android_external_format_resolve_spec_version = 1
pub const android_external_format_resolve_extension_name = "VK_ANDROID_external_format_resolve"
// PhysicalDeviceExternalFormatResolveFeaturesANDROID extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceExternalFormatResolveFeaturesANDROID {
mut:
    s_type                 StructureType
    p_next                 voidptr
    external_format_resolve Bool32
} 

// PhysicalDeviceExternalFormatResolvePropertiesANDROID extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceExternalFormatResolvePropertiesANDROID {
mut:
    s_type                  StructureType
    p_next                  voidptr
    null_color_attachment_with_external_format_resolve Bool32
    external_format_resolve_chroma_offset_x ChromaLocation
    external_format_resolve_chroma_offset_y ChromaLocation
} 

// AndroidHardwareBufferFormatResolvePropertiesANDROID extends VkAndroidHardwareBufferPropertiesANDROID
pub struct AndroidHardwareBufferFormatResolvePropertiesANDROID {
mut:
    s_type                 StructureType
    p_next                 voidptr
    color_attachment_format Format
} 



// VK_EXT_shader_object is a preprocessor guard. Do not pass it to API calls.
const ext_shader_object = 1
pub type C.ShaderEXT = voidptr
pub const ext_shader_object_spec_version    = 1
pub const ext_shader_object_extension_name  = "VK_EXT_shader_object"

pub enum ShaderCodeTypeEXT {
    shader_code_type_binary_ext = int(0)
    shader_code_type_spirv_ext = int(1)
    shader_code_type_max_enum_ext = int(0x7FFFFFFF)
}


pub enum ShaderCreateFlagBitsEXT {
    shader_create_link_stage_bit_ext = int(0x00000001)
    shader_create_allow_varying_subgroup_size_bit_ext = int(0x00000002)
    shader_create_require_full_subgroups_bit_ext = int(0x00000004)
    shader_create_no_task_shader_bit_ext = int(0x00000008)
    shader_create_dispatch_base_bit_ext = int(0x00000010)
    shader_create_fragment_shading_rate_attachment_bit_ext = int(0x00000020)
    shader_create_fragment_density_map_attachment_bit_ext = int(0x00000040)
    shader_create_flag_bits_max_enum_ext = int(0x7FFFFFFF)
}

pub type ShaderCreateFlagsEXT = u32
// PhysicalDeviceShaderObjectFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderObjectFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_object          Bool32
} 

// PhysicalDeviceShaderObjectPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceShaderObjectPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_binary_uuid     []u8
    shader_binary_version  u32
} 

pub struct ShaderCreateInfoEXT {
mut:
    s_type                              StructureType
    p_next                              voidptr
    flags                               ShaderCreateFlagsEXT
    stage                               ShaderStageFlagBits
    next_stage                          ShaderStageFlags
    code_type                           ShaderCodeTypeEXT
    code_size                           usize
    p_code                              voidptr
    p_name                              &char
    set_layout_count                    u32
    p_set_layouts                       &C.DescriptorSetLayout
    push_constant_range_count           u32
    p_push_constant_ranges              &PushConstantRange
    p_specialization_info               &SpecializationInfo
} 

pub type ShaderRequiredSubgroupSizeCreateInfoEXT = PipelineShaderStageRequiredSubgroupSizeCreateInfo

type VkCreateShadersEXT = fn (     C.Device,     u32,     &ShaderCreateInfoEXT,     &AllocationCallbacks,     &C.ShaderEXT) Result

pub fn create_shaders_ext(
    device                                          C.Device,
    create_info_count                               u32,
    p_create_infos                                  &ShaderCreateInfoEXT,
    p_allocator                                     &AllocationCallbacks,
    p_shaders                                       &C.ShaderEXT) Result {
      f := VkCreateShadersEXT((*loader_p).get_sym('vkCreateShadersEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCreateShadersEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    create_info_count,
    p_create_infos,
    p_allocator,
    p_shaders)
}


type VkDestroyShaderEXT = fn (     C.Device,     C.ShaderEXT,     &AllocationCallbacks) 

pub fn destroy_shader_ext(
    device                                          C.Device,
    shader                                          C.ShaderEXT,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyShaderEXT((*loader_p).get_sym('vkDestroyShaderEXT'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyShaderEXT': ${err}")
        return 
    })
    f(
    device,
    shader,
    p_allocator)
}


type VkGetShaderBinaryDataEXT = fn (     C.Device,     C.ShaderEXT,     &usize,     voidptr) Result

pub fn get_shader_binary_data_ext(
    device                                          C.Device,
    shader                                          C.ShaderEXT,
    p_data_size                                     &usize,
    p_data                                          voidptr) Result {
      f := VkGetShaderBinaryDataEXT((*loader_p).get_sym('vkGetShaderBinaryDataEXT'
    ) or { 
        println("Couldn't load symbol for 'vkGetShaderBinaryDataEXT': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    shader,
    p_data_size,
    p_data)
}


type VkCmdBindShadersEXT = fn (     C.CommandBuffer,     u32,     &ShaderStageFlagBits,     &C.ShaderEXT) 

pub fn cmd_bind_shaders_ext(
    command_buffer                                  C.CommandBuffer,
    stage_count                                     u32,
    p_stages                                        &ShaderStageFlagBits,
    p_shaders                                       &C.ShaderEXT)  {
      f := VkCmdBindShadersEXT((*loader_p).get_sym('vkCmdBindShadersEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBindShadersEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    stage_count,
    p_stages,
    p_shaders)
}




// VK_QCOM_tile_properties is a preprocessor guard. Do not pass it to API calls.
const qcom_tile_properties = 1
pub const qcom_tile_properties_spec_version = 1
pub const qcom_tile_properties_extension_name = "VK_QCOM_tile_properties"
// PhysicalDeviceTilePropertiesFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceTilePropertiesFeaturesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    tile_properties        Bool32
} 

pub struct TilePropertiesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    tile_size              Extent3D
    apron_size             Extent2D
    origin                 Offset2D
} 

type VkGetFramebufferTilePropertiesQCOM = fn (     C.Device,     C.Framebuffer,     &u32,     &TilePropertiesQCOM) Result

pub fn get_framebuffer_tile_properties_qcom(
    device                                          C.Device,
    framebuffer                                     C.Framebuffer,
    p_properties_count                              &u32,
    p_properties                                    &TilePropertiesQCOM) Result {
      f := VkGetFramebufferTilePropertiesQCOM((*loader_p).get_sym('vkGetFramebufferTilePropertiesQCOM'
    ) or { 
        println("Couldn't load symbol for 'vkGetFramebufferTilePropertiesQCOM': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    framebuffer,
    p_properties_count,
    p_properties)
}


type VkGetDynamicRenderingTilePropertiesQCOM = fn (     C.Device,     &RenderingInfo,     &TilePropertiesQCOM) Result

pub fn get_dynamic_rendering_tile_properties_qcom(
    device                                          C.Device,
    p_rendering_info                                &RenderingInfo,
    p_properties                                    &TilePropertiesQCOM) Result {
      f := VkGetDynamicRenderingTilePropertiesQCOM((*loader_p).get_sym('vkGetDynamicRenderingTilePropertiesQCOM'
    ) or { 
        println("Couldn't load symbol for 'vkGetDynamicRenderingTilePropertiesQCOM': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_rendering_info,
    p_properties)
}




// VK_SEC_amigo_profiling is a preprocessor guard. Do not pass it to API calls.
const sec_amigo_profiling = 1
pub const sec_amigo_profiling_spec_version  = 1
pub const sec_amigo_profiling_extension_name = "VK_SEC_amigo_profiling"
// PhysicalDeviceAmigoProfilingFeaturesSEC extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceAmigoProfilingFeaturesSEC {
mut:
    s_type                 StructureType
    p_next                 voidptr
    amigo_profiling        Bool32
} 

// AmigoProfilingSubmitInfoSEC extends VkSubmitInfo
pub struct AmigoProfilingSubmitInfoSEC {
mut:
    s_type                 StructureType
    p_next                 voidptr
    first_draw_timestamp   u64
    swap_buffer_timestamp  u64
} 



// VK_QCOM_multiview_per_view_viewports is a preprocessor guard. Do not pass it to API calls.
const qcom_multiview_per_view_viewports = 1
pub const qcom_multiview_per_view_viewports_spec_version = 1
pub const qcom_multiview_per_view_viewports_extension_name = "VK_QCOM_multiview_per_view_viewports"
// PhysicalDeviceMultiviewPerViewViewportsFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMultiviewPerViewViewportsFeaturesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    multiview_per_view_viewports Bool32
} 



// VK_NV_ray_tracing_invocation_reorder is a preprocessor guard. Do not pass it to API calls.
const nv_ray_tracing_invocation_reorder = 1
pub const nv_ray_tracing_invocation_reorder_spec_version = 1
pub const nv_ray_tracing_invocation_reorder_extension_name = "VK_NV_ray_tracing_invocation_reorder"

pub enum RayTracingInvocationReorderModeNV {
    ray_tracing_invocation_reorder_mode_none_nv = int(0)
    ray_tracing_invocation_reorder_mode_reorder_nv = int(1)
    ray_tracing_invocation_reorder_mode_max_enum_nv = int(0x7FFFFFFF)
}

// PhysicalDeviceRayTracingInvocationReorderPropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceRayTracingInvocationReorderPropertiesNV {
mut:
    s_type                                     StructureType
    p_next                                     voidptr
    ray_tracing_invocation_reorder_reordering_hint RayTracingInvocationReorderModeNV
} 

// PhysicalDeviceRayTracingInvocationReorderFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRayTracingInvocationReorderFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    ray_tracing_invocation_reorder Bool32
} 



// VK_NV_extended_sparse_address_space is a preprocessor guard. Do not pass it to API calls.
const nv_extended_sparse_address_space = 1
pub const nv_extended_sparse_address_space_spec_version = 1
pub const nv_extended_sparse_address_space_extension_name = "VK_NV_extended_sparse_address_space"
// PhysicalDeviceExtendedSparseAddressSpaceFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceExtendedSparseAddressSpaceFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    extended_sparse_address_space Bool32
} 

// PhysicalDeviceExtendedSparseAddressSpacePropertiesNV extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceExtendedSparseAddressSpacePropertiesNV {
mut:
    s_type                    StructureType
    p_next                    voidptr
    extended_sparse_address_space_size DeviceSize
    extended_sparse_image_usage_flags ImageUsageFlags
    extended_sparse_buffer_usage_flags BufferUsageFlags
} 



// VK_EXT_mutable_descriptor_type is a preprocessor guard. Do not pass it to API calls.
const ext_mutable_descriptor_type = 1
pub const ext_mutable_descriptor_type_spec_version = 1
pub const ext_mutable_descriptor_type_extension_name = "VK_EXT_mutable_descriptor_type"


// VK_EXT_layer_settings is a preprocessor guard. Do not pass it to API calls.
const ext_layer_settings = 1
pub const ext_layer_settings_spec_version   = 2
pub const ext_layer_settings_extension_name = "VK_EXT_layer_settings"

pub enum LayerSettingTypeEXT {
    layer_setting_type_bool32_ext = int(0)
    layer_setting_type_int32_ext = int(1)
    layer_setting_type_int64_ext = int(2)
    layer_setting_type_uint32_ext = int(3)
    layer_setting_type_uint64_ext = int(4)
    layer_setting_type_float32_ext = int(5)
    layer_setting_type_float64_ext = int(6)
    layer_setting_type_string_ext = int(7)
    layer_setting_type_max_enum_ext = int(0x7FFFFFFF)
}

pub struct LayerSettingEXT {
mut:
    p_layer_name                 &char
    p_setting_name               &char
    vktype                       LayerSettingTypeEXT
    value_count                  u32
    p_values                     voidptr
} 

// LayerSettingsCreateInfoEXT extends VkInstanceCreateInfo
pub struct LayerSettingsCreateInfoEXT {
mut:
    s_type                          StructureType
    p_next                          voidptr
    setting_count                   u32
    p_settings                      &LayerSettingEXT
} 



// VK_ARM_shader_core_builtins is a preprocessor guard. Do not pass it to API calls.
const arm_shader_core_builtins = 1
pub const arm_shader_core_builtins_spec_version = 2
pub const arm_shader_core_builtins_extension_name = "VK_ARM_shader_core_builtins"
// PhysicalDeviceShaderCoreBuiltinsFeaturesARM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceShaderCoreBuiltinsFeaturesARM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_core_builtins   Bool32
} 

// PhysicalDeviceShaderCoreBuiltinsPropertiesARM extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceShaderCoreBuiltinsPropertiesARM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_core_mask       u64
    shader_core_count      u32
    shader_warps_per_core  u32
} 



// VK_EXT_pipeline_library_group_handles is a preprocessor guard. Do not pass it to API calls.
const ext_pipeline_library_group_handles = 1
pub const ext_pipeline_library_group_handles_spec_version = 1
pub const ext_pipeline_library_group_handles_extension_name = "VK_EXT_pipeline_library_group_handles"
// PhysicalDevicePipelineLibraryGroupHandlesFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDevicePipelineLibraryGroupHandlesFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    pipeline_library_group_handles Bool32
} 



// VK_EXT_dynamic_rendering_unused_attachments is a preprocessor guard. Do not pass it to API calls.
const ext_dynamic_rendering_unused_attachments = 1
pub const ext_dynamic_rendering_unused_attachments_spec_version = 1
pub const ext_dynamic_rendering_unused_attachments_extension_name = "VK_EXT_dynamic_rendering_unused_attachments"
// PhysicalDeviceDynamicRenderingUnusedAttachmentsFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDynamicRenderingUnusedAttachmentsFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    dynamic_rendering_unused_attachments Bool32
} 



// VK_NV_low_latency2 is a preprocessor guard. Do not pass it to API calls.
const nv_low_latency2 = 1
pub const nv_low_latency_2_spec_version     = 2
pub const nv_low_latency_2_extension_name   = "VK_NV_low_latency2"

pub enum LatencyMarkerNV {
    latency_marker_simulation_start_nv = int(0)
    latency_marker_simulation_end_nv = int(1)
    latency_marker_rendersubmit_start_nv = int(2)
    latency_marker_rendersubmit_end_nv = int(3)
    latency_marker_present_start_nv = int(4)
    latency_marker_present_end_nv = int(5)
    latency_marker_input_sample_nv = int(6)
    latency_marker_trigger_flash_nv = int(7)
    latency_marker_out_of_band_rendersubmit_start_nv = int(8)
    latency_marker_out_of_band_rendersubmit_end_nv = int(9)
    latency_marker_out_of_band_present_start_nv = int(10)
    latency_marker_out_of_band_present_end_nv = int(11)
    latency_marker_max_enum_nv = int(0x7FFFFFFF)
}


pub enum OutOfBandQueueTypeNV {
    out_of_band_queue_type_render_nv = int(0)
    out_of_band_queue_type_present_nv = int(1)
    out_of_band_queue_type_max_enum_nv = int(0x7FFFFFFF)
}

pub struct LatencySleepModeInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    low_latency_mode       Bool32
    low_latency_boost      Bool32
    minimum_interval_us    u32
} 

pub struct LatencySleepInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    signal_semaphore       C.Semaphore
    value                  u64
} 

pub struct SetLatencyMarkerInfoNV {
mut:
    s_type                   StructureType
    p_next                   voidptr
    present_id               u64
    marker                   LatencyMarkerNV
} 

pub struct LatencyTimingsFrameReportNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    present_id             u64
    input_sample_time_us   u64
    sim_start_time_us      u64
    sim_end_time_us        u64
    render_submit_start_time_us u64
    render_submit_end_time_us u64
    present_start_time_us  u64
    present_end_time_us    u64
    driver_start_time_us   u64
    driver_end_time_us     u64
    os_render_queue_start_time_us u64
    os_render_queue_end_time_us u64
    gpu_render_start_time_us u64
    gpu_render_end_time_us u64
} 

pub struct GetLatencyMarkerInfoNV {
mut:
    s_type                                StructureType
    p_next                                voidptr
    timing_count                          u32
    p_timings                             &LatencyTimingsFrameReportNV
} 

// LatencySubmissionPresentIdNV extends VkSubmitInfo,VkSubmitInfo2
pub struct LatencySubmissionPresentIdNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    present_id             u64
} 

// SwapchainLatencyCreateInfoNV extends VkSwapchainCreateInfoKHR
pub struct SwapchainLatencyCreateInfoNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    latency_mode_enable    Bool32
} 

pub struct OutOfBandQueueTypeInfoNV {
mut:
    s_type                        StructureType
    p_next                        voidptr
    queue_type                    OutOfBandQueueTypeNV
} 

// LatencySurfaceCapabilitiesNV extends VkSurfaceCapabilities2KHR
pub struct LatencySurfaceCapabilitiesNV {
mut:
    s_type                   StructureType
    p_next                   voidptr
    present_mode_count       u32
    p_present_modes          &PresentModeKHR
} 

type VkSetLatencySleepModeNV = fn (     C.Device,     C.SwapchainKHR,     &LatencySleepModeInfoNV) Result

pub fn set_latency_sleep_mode_nv(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR,
    p_sleep_mode_info                               &LatencySleepModeInfoNV) Result {
      f := VkSetLatencySleepModeNV((*loader_p).get_sym('vkSetLatencySleepModeNV'
    ) or { 
        println("Couldn't load symbol for 'vkSetLatencySleepModeNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain,
    p_sleep_mode_info)
}


type VkLatencySleepNV = fn (     C.Device,     C.SwapchainKHR,     &LatencySleepInfoNV) Result

pub fn latency_sleep_nv(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR,
    p_sleep_info                                    &LatencySleepInfoNV) Result {
      f := VkLatencySleepNV((*loader_p).get_sym('vkLatencySleepNV'
    ) or { 
        println("Couldn't load symbol for 'vkLatencySleepNV': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    swapchain,
    p_sleep_info)
}


type VkSetLatencyMarkerNV = fn (     C.Device,     C.SwapchainKHR,     &SetLatencyMarkerInfoNV) 

pub fn set_latency_marker_nv(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR,
    p_latency_marker_info                           &SetLatencyMarkerInfoNV)  {
      f := VkSetLatencyMarkerNV((*loader_p).get_sym('vkSetLatencyMarkerNV'
    ) or { 
        println("Couldn't load symbol for 'vkSetLatencyMarkerNV': ${err}")
        return 
    })
    f(
    device,
    swapchain,
    p_latency_marker_info)
}


type VkGetLatencyTimingsNV = fn (     C.Device,     C.SwapchainKHR,     &GetLatencyMarkerInfoNV) 

pub fn get_latency_timings_nv(
    device                                          C.Device,
    swapchain                                       C.SwapchainKHR,
    p_latency_marker_info                           &GetLatencyMarkerInfoNV)  {
      f := VkGetLatencyTimingsNV((*loader_p).get_sym('vkGetLatencyTimingsNV'
    ) or { 
        println("Couldn't load symbol for 'vkGetLatencyTimingsNV': ${err}")
        return 
    })
    f(
    device,
    swapchain,
    p_latency_marker_info)
}


type VkQueueNotifyOutOfBandNV = fn (     C.Queue,     &OutOfBandQueueTypeInfoNV) 

pub fn queue_notify_out_of_band_nv(
    queue                                           C.Queue,
    p_queue_type_info                               &OutOfBandQueueTypeInfoNV)  {
      f := VkQueueNotifyOutOfBandNV((*loader_p).get_sym('vkQueueNotifyOutOfBandNV'
    ) or { 
        println("Couldn't load symbol for 'vkQueueNotifyOutOfBandNV': ${err}")
        return 
    })
    f(
    queue,
    p_queue_type_info)
}




// VK_QCOM_multiview_per_view_render_areas is a preprocessor guard. Do not pass it to API calls.
const qcom_multiview_per_view_render_areas = 1
pub const qcom_multiview_per_view_render_areas_spec_version = 1
pub const qcom_multiview_per_view_render_areas_extension_name = "VK_QCOM_multiview_per_view_render_areas"
// PhysicalDeviceMultiviewPerViewRenderAreasFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMultiviewPerViewRenderAreasFeaturesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    multiview_per_view_render_areas Bool32
} 

// MultiviewPerViewRenderAreasRenderPassBeginInfoQCOM extends VkRenderPassBeginInfo,VkRenderingInfo
pub struct MultiviewPerViewRenderAreasRenderPassBeginInfoQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    per_view_render_area_count u32
    p_per_view_render_areas &Rect2D
} 



// VK_QCOM_image_processing2 is a preprocessor guard. Do not pass it to API calls.
const qcom_image_processing2 = 1
pub const qcom_image_processing_2_spec_version = 1
pub const qcom_image_processing_2_extension_name = "VK_QCOM_image_processing2"

pub enum BlockMatchWindowCompareModeQCOM {
    block_match_window_compare_mode_min_qcom = int(0)
    block_match_window_compare_mode_max_qcom = int(1)
    block_match_window_compare_mode_max_enum_qcom = int(0x7FFFFFFF)
}

// PhysicalDeviceImageProcessing2FeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceImageProcessing2FeaturesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    texture_block_match2   Bool32
} 

// PhysicalDeviceImageProcessing2PropertiesQCOM extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceImageProcessing2PropertiesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_block_match_window Extent2D
} 

// SamplerBlockMatchWindowCreateInfoQCOM extends VkSamplerCreateInfo
pub struct SamplerBlockMatchWindowCreateInfoQCOM {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    window_extent                            Extent2D
    window_compare_mode                      BlockMatchWindowCompareModeQCOM
} 



// VK_QCOM_filter_cubic_weights is a preprocessor guard. Do not pass it to API calls.
const qcom_filter_cubic_weights = 1
pub const qcom_filter_cubic_weights_spec_version = 1
pub const qcom_filter_cubic_weights_extension_name = "VK_QCOM_filter_cubic_weights"

pub enum CubicFilterWeightsQCOM {
    cubic_filter_weights_catmull_rom_qcom = int(0)
    cubic_filter_weights_zero_tangent_cardinal_qcom = int(1)
    cubic_filter_weights_b_spline_qcom = int(2)
    cubic_filter_weights_mitchell_netravali_qcom = int(3)
    cubic_filter_weights_max_enum_qcom = int(0x7FFFFFFF)
}

// PhysicalDeviceCubicWeightsFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceCubicWeightsFeaturesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    selectable_cubic_weights Bool32
} 

// SamplerCubicWeightsCreateInfoQCOM extends VkSamplerCreateInfo
pub struct SamplerCubicWeightsCreateInfoQCOM {
mut:
    s_type                          StructureType
    p_next                          voidptr
    cubic_weights                   CubicFilterWeightsQCOM
} 

// BlitImageCubicWeightsInfoQCOM extends VkBlitImageInfo2
pub struct BlitImageCubicWeightsInfoQCOM {
mut:
    s_type                          StructureType
    p_next                          voidptr
    cubic_weights                   CubicFilterWeightsQCOM
} 



// VK_QCOM_ycbcr_degamma is a preprocessor guard. Do not pass it to API calls.
const qcom_ycbcr_degamma = 1
pub const qcom_ycbcr_degamma_spec_version   = 1
pub const qcom_ycbcr_degamma_extension_name = "VK_QCOM_ycbcr_degamma"
// PhysicalDeviceYcbcrDegammaFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceYcbcrDegammaFeaturesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    ycbcr_degamma          Bool32
} 

// SamplerYcbcrConversionYcbcrDegammaCreateInfoQCOM extends VkSamplerYcbcrConversionCreateInfo
pub struct SamplerYcbcrConversionYcbcrDegammaCreateInfoQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    enable_y_degamma       Bool32
    enable_cb_cr_degamma   Bool32
} 



// VK_QCOM_filter_cubic_clamp is a preprocessor guard. Do not pass it to API calls.
const qcom_filter_cubic_clamp = 1
pub const qcom_filter_cubic_clamp_spec_version = 1
pub const qcom_filter_cubic_clamp_extension_name = "VK_QCOM_filter_cubic_clamp"
// PhysicalDeviceCubicClampFeaturesQCOM extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceCubicClampFeaturesQCOM {
mut:
    s_type                 StructureType
    p_next                 voidptr
    cubic_range_clamp      Bool32
} 



// VK_EXT_attachment_feedback_loop_dynamic_state is a preprocessor guard. Do not pass it to API calls.
const ext_attachment_feedback_loop_dynamic_state = 1
pub const ext_attachment_feedback_loop_dynamic_state_spec_version = 1
pub const ext_attachment_feedback_loop_dynamic_state_extension_name = "VK_EXT_attachment_feedback_loop_dynamic_state"
// PhysicalDeviceAttachmentFeedbackLoopDynamicStateFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceAttachmentFeedbackLoopDynamicStateFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    attachment_feedback_loop_dynamic_state Bool32
} 

type VkCmdSetAttachmentFeedbackLoopEnableEXT = fn (     C.CommandBuffer,     ImageAspectFlags) 

pub fn cmd_set_attachment_feedback_loop_enable_ext(
    command_buffer                                  C.CommandBuffer,
    aspect_mask                                     ImageAspectFlags)  {
      f := VkCmdSetAttachmentFeedbackLoopEnableEXT((*loader_p).get_sym('vkCmdSetAttachmentFeedbackLoopEnableEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetAttachmentFeedbackLoopEnableEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    aspect_mask)
}




// VK_QNX_external_memory_screen_buffer is a preprocessor guard. Do not pass it to API calls.
const qnx_external_memory_screen_buffer = 1
pub const qnx_external_memory_screen_buffer_spec_version = 1
pub const qnx_external_memory_screen_buffer_extension_name = "VK_QNX_external_memory_screen_buffer"
pub struct ScreenBufferPropertiesQNX {
mut:
    s_type                 StructureType
    p_next                 voidptr
    allocation_size        DeviceSize
    memory_type_bits       u32
} 

// ScreenBufferFormatPropertiesQNX extends VkScreenBufferPropertiesQNX
pub struct ScreenBufferFormatPropertiesQNX {
mut:
    s_type                               StructureType
    p_next                               voidptr
    format                               Format
    external_format                      u64
    screen_usage                         u64
    format_features                      FormatFeatureFlags
    sampler_ycbcr_conversion_components  ComponentMapping
    suggested_ycbcr_model                SamplerYcbcrModelConversion
    suggested_ycbcr_range                SamplerYcbcrRange
    suggested_x_chroma_offset            ChromaLocation
    suggested_y_chroma_offset            ChromaLocation
} 

// ImportScreenBufferInfoQNX extends VkMemoryAllocateInfo
pub struct ImportScreenBufferInfoQNX {
mut:
    s_type                        StructureType
    p_next                        voidptr
    buffer                        voidptr
} 

// ExternalFormatQNX extends VkImageCreateInfo,VkSamplerYcbcrConversionCreateInfo
pub struct ExternalFormatQNX {
mut:
    s_type                 StructureType
    p_next                 voidptr
    external_format        u64
} 

// PhysicalDeviceExternalMemoryScreenBufferFeaturesQNX extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceExternalMemoryScreenBufferFeaturesQNX {
mut:
    s_type                 StructureType
    p_next                 voidptr
    screen_buffer_import   Bool32
} 

type VkGetScreenBufferPropertiesQNX = fn (     C.Device,     voidptr,     &ScreenBufferPropertiesQNX) Result

pub fn get_screen_buffer_properties_qnx(
    device                                          C.Device,
    buffer                                          voidptr,
    p_properties                                    &ScreenBufferPropertiesQNX) Result {
      f := VkGetScreenBufferPropertiesQNX((*loader_p).get_sym('vkGetScreenBufferPropertiesQNX'
    ) or { 
        println("Couldn't load symbol for 'vkGetScreenBufferPropertiesQNX': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    buffer,
    p_properties)
}




// VK_MSFT_layered_driver is a preprocessor guard. Do not pass it to API calls.
const msft_layered_driver = 1
pub const msft_layered_driver_spec_version  = 1
pub const msft_layered_driver_extension_name = "VK_MST_layered_driver"

pub enum LayeredDriverUnderlyingApiMSFT {
    layered_driver_underlying_api_none_msft = int(0)
    layered_driver_underlying_api_d3d12_msft = int(1)
    layered_driver_underlying_api_max_enum_msft = int(0x7FFFFFFF)
}

// PhysicalDeviceLayeredDriverPropertiesMSFT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceLayeredDriverPropertiesMSFT {
mut:
    s_type                                  StructureType
    p_next                                  voidptr
    underlying_api                          LayeredDriverUnderlyingApiMSFT
} 



// VK_NV_descriptor_pool_overallocation is a preprocessor guard. Do not pass it to API calls.
const nv_descriptor_pool_overallocation = 1
pub const nv_descriptor_pool_overallocation_spec_version = 1
pub const nv_descriptor_pool_overallocation_extension_name = "VK_NV_descriptor_pool_overallocation"
// PhysicalDeviceDescriptorPoolOverallocationFeaturesNV extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceDescriptorPoolOverallocationFeaturesNV {
mut:
    s_type                 StructureType
    p_next                 voidptr
    descriptor_pool_overallocation Bool32
} 



// VK_KHR_acceleration_structure is a preprocessor guard. Do not pass it to API calls.
const khr_acceleration_structure = 1
pub const khr_acceleration_structure_spec_version = 13
pub const khr_acceleration_structure_extension_name = "VK_KHR_acceleration_structure"

pub enum BuildAccelerationStructureModeKHR {
    build_acceleration_structure_mode_build_khr = int(0)
    build_acceleration_structure_mode_update_khr = int(1)
    build_acceleration_structure_mode_max_enum_khr = int(0x7FFFFFFF)
}


pub enum AccelerationStructureCreateFlagBitsKHR {
    acceleration_structure_create_device_address_capture_replay_bit_khr = int(0x00000001)
    acceleration_structure_create_descriptor_buffer_capture_replay_bit_ext = int(0x00000008)
    acceleration_structure_create_motion_bit_nv = int(0x00000004)
    acceleration_structure_create_flag_bits_max_enum_khr = int(0x7FFFFFFF)
}

pub type AccelerationStructureCreateFlagsKHR = u32
pub struct AccelerationStructureBuildRangeInfoKHR {
mut:
    primitive_count u32
    primitive_offset u32
    first_vertex    u32
    transform_offset u32
} 

pub struct AccelerationStructureGeometryTrianglesDataKHR {
mut:
    s_type                               StructureType
    p_next                               voidptr
    vertex_format                        Format
    vertex_data                          DeviceOrHostAddressConstKHR
    vertex_stride                        DeviceSize
    max_vertex                           u32
    index_type                           IndexType
    index_data                           DeviceOrHostAddressConstKHR
    transform_data                       DeviceOrHostAddressConstKHR
} 

pub struct AccelerationStructureGeometryAabbsDataKHR {
mut:
    s_type                               StructureType
    p_next                               voidptr
    data                                 DeviceOrHostAddressConstKHR
    stride                               DeviceSize
} 

pub struct AccelerationStructureGeometryInstancesDataKHR {
mut:
    s_type                               StructureType
    p_next                               voidptr
    array_of_pointers                    Bool32
    data                                 DeviceOrHostAddressConstKHR
} 

pub union AccelerationStructureGeometryDataKHR {
mut:
    triangles                                              AccelerationStructureGeometryTrianglesDataKHR
    aabbs                                                  AccelerationStructureGeometryAabbsDataKHR
    instances                                              AccelerationStructureGeometryInstancesDataKHR
} 

pub struct AccelerationStructureGeometryKHR {
mut:
    s_type                                        StructureType
    p_next                                        voidptr
    geometry_type                                 GeometryTypeKHR
    geometry                                      AccelerationStructureGeometryDataKHR
    flags                                         GeometryFlagsKHR
} 

pub struct AccelerationStructureBuildGeometryInfoKHR {
mut:
    s_type                                                  StructureType
    p_next                                                  voidptr
    vktype                                                  AccelerationStructureTypeKHR
    flags                                                   BuildAccelerationStructureFlagsKHR
    mode                                                    BuildAccelerationStructureModeKHR
    src_acceleration_structure                              C.AccelerationStructureKHR
    dst_acceleration_structure                              C.AccelerationStructureKHR
    geometry_count                                          u32
    p_geometries                                            &AccelerationStructureGeometryKHR
    pp_geometries                                           &AccelerationStructureGeometryKHR
    scratch_data                                            DeviceOrHostAddressKHR
} 

pub struct AccelerationStructureCreateInfoKHR {
mut:
    s_type                                       StructureType
    p_next                                       voidptr
    create_flags                                 AccelerationStructureCreateFlagsKHR
    buffer                                       C.Buffer
    offset                                       DeviceSize
    size                                         DeviceSize
    vktype                                       AccelerationStructureTypeKHR
    device_address                               DeviceAddress
} 

// WriteDescriptorSetAccelerationStructureKHR extends VkWriteDescriptorSet
pub struct WriteDescriptorSetAccelerationStructureKHR {
mut:
    s_type                                   StructureType
    p_next                                   voidptr
    acceleration_structure_count             u32
    p_acceleration_structures                &C.AccelerationStructureKHR
} 

// PhysicalDeviceAccelerationStructureFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceAccelerationStructureFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    acceleration_structure Bool32
    acceleration_structure_capture_replay Bool32
    acceleration_structure_indirect_build Bool32
    acceleration_structure_host_commands Bool32
    descriptor_binding_acceleration_structure_update_after_bind Bool32
} 

// PhysicalDeviceAccelerationStructurePropertiesKHR extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceAccelerationStructurePropertiesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_geometry_count     u64
    max_instance_count     u64
    max_primitive_count    u64
    max_per_stage_descriptor_acceleration_structures u32
    max_per_stage_descriptor_update_after_bind_acceleration_structures u32
    max_descriptor_set_acceleration_structures u32
    max_descriptor_set_update_after_bind_acceleration_structures u32
    min_acceleration_structure_scratch_offset_alignment u32
} 

pub struct AccelerationStructureDeviceAddressInfoKHR {
mut:
    s_type                            StructureType
    p_next                            voidptr
    acceleration_structure            C.AccelerationStructureKHR
} 

pub struct AccelerationStructureVersionInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    p_version_data         &u8
} 

pub struct CopyAccelerationStructureToMemoryInfoKHR {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    src                                       C.AccelerationStructureKHR
    dst                                       DeviceOrHostAddressKHR
    mode                                      CopyAccelerationStructureModeKHR
} 

pub struct CopyMemoryToAccelerationStructureInfoKHR {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    src                                       DeviceOrHostAddressConstKHR
    dst                                       C.AccelerationStructureKHR
    mode                                      CopyAccelerationStructureModeKHR
} 

pub struct CopyAccelerationStructureInfoKHR {
mut:
    s_type                                    StructureType
    p_next                                    voidptr
    src                                       C.AccelerationStructureKHR
    dst                                       C.AccelerationStructureKHR
    mode                                      CopyAccelerationStructureModeKHR
} 

pub struct AccelerationStructureBuildSizesInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    acceleration_structure_size DeviceSize
    update_scratch_size    DeviceSize
    build_scratch_size     DeviceSize
} 

type VkCreateAccelerationStructureKHR = fn (     C.Device,     &AccelerationStructureCreateInfoKHR,     &AllocationCallbacks,     &C.AccelerationStructureKHR) Result

pub fn create_acceleration_structure_khr(
    device                                          C.Device,
    p_create_info                                   &AccelerationStructureCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_acceleration_structure                        &C.AccelerationStructureKHR) Result {
      f := VkCreateAccelerationStructureKHR((*loader_p).get_sym('vkCreateAccelerationStructureKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateAccelerationStructureKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    p_create_info,
    p_allocator,
    p_acceleration_structure)
}


type VkDestroyAccelerationStructureKHR = fn (     C.Device,     C.AccelerationStructureKHR,     &AllocationCallbacks) 

pub fn destroy_acceleration_structure_khr(
    device                                          C.Device,
    acceleration_structure                          C.AccelerationStructureKHR,
    p_allocator                                     &AllocationCallbacks)  {
      f := VkDestroyAccelerationStructureKHR((*loader_p).get_sym('vkDestroyAccelerationStructureKHR'
    ) or { 
        println("Couldn't load symbol for 'vkDestroyAccelerationStructureKHR': ${err}")
        return 
    })
    f(
    device,
    acceleration_structure,
    p_allocator)
}


type VkCmdBuildAccelerationStructuresKHR = fn (     C.CommandBuffer,     u32,     &AccelerationStructureBuildGeometryInfoKHR,     &AccelerationStructureBuildRangeInfoKHR) 

pub fn cmd_build_acceleration_structures_khr(
    command_buffer                                  C.CommandBuffer,
    info_count                                      u32,
    p_infos                                         &AccelerationStructureBuildGeometryInfoKHR,
    pp_build_range_infos                            &AccelerationStructureBuildRangeInfoKHR)  {
      f := VkCmdBuildAccelerationStructuresKHR((*loader_p).get_sym('vkCmdBuildAccelerationStructuresKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBuildAccelerationStructuresKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    info_count,
    p_infos,
    pp_build_range_infos)
}


type VkCmdBuildAccelerationStructuresIndirectKHR = fn (     C.CommandBuffer,     u32,     &AccelerationStructureBuildGeometryInfoKHR,     &DeviceAddress,     &u32,     &u32) 

pub fn cmd_build_acceleration_structures_indirect_khr(
    command_buffer                                  C.CommandBuffer,
    info_count                                      u32,
    p_infos                                         &AccelerationStructureBuildGeometryInfoKHR,
    p_indirect_device_addresses                     &DeviceAddress,
    p_indirect_strides                              &u32,
    pp_max_primitive_counts                         &u32)  {
      f := VkCmdBuildAccelerationStructuresIndirectKHR((*loader_p).get_sym('vkCmdBuildAccelerationStructuresIndirectKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdBuildAccelerationStructuresIndirectKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    info_count,
    p_infos,
    p_indirect_device_addresses,
    p_indirect_strides,
    pp_max_primitive_counts)
}


type VkBuildAccelerationStructuresKHR = fn (     C.Device,     C.DeferredOperationKHR,     u32,     &AccelerationStructureBuildGeometryInfoKHR,     &AccelerationStructureBuildRangeInfoKHR) Result

pub fn build_acceleration_structures_khr(
    device                                          C.Device,
    deferred_operation                              C.DeferredOperationKHR,
    info_count                                      u32,
    p_infos                                         &AccelerationStructureBuildGeometryInfoKHR,
    pp_build_range_infos                            &AccelerationStructureBuildRangeInfoKHR) Result {
      f := VkBuildAccelerationStructuresKHR((*loader_p).get_sym('vkBuildAccelerationStructuresKHR'
    ) or { 
        println("Couldn't load symbol for 'vkBuildAccelerationStructuresKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    deferred_operation,
    info_count,
    p_infos,
    pp_build_range_infos)
}


type VkCopyAccelerationStructureKHR = fn (     C.Device,     C.DeferredOperationKHR,     &CopyAccelerationStructureInfoKHR) Result

pub fn copy_acceleration_structure_khr(
    device                                          C.Device,
    deferred_operation                              C.DeferredOperationKHR,
    p_info                                          &CopyAccelerationStructureInfoKHR) Result {
      f := VkCopyAccelerationStructureKHR((*loader_p).get_sym('vkCopyAccelerationStructureKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCopyAccelerationStructureKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    deferred_operation,
    p_info)
}


type VkCopyAccelerationStructureToMemoryKHR = fn (     C.Device,     C.DeferredOperationKHR,     &CopyAccelerationStructureToMemoryInfoKHR) Result

pub fn copy_acceleration_structure_to_memory_khr(
    device                                          C.Device,
    deferred_operation                              C.DeferredOperationKHR,
    p_info                                          &CopyAccelerationStructureToMemoryInfoKHR) Result {
      f := VkCopyAccelerationStructureToMemoryKHR((*loader_p).get_sym('vkCopyAccelerationStructureToMemoryKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCopyAccelerationStructureToMemoryKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    deferred_operation,
    p_info)
}


type VkCopyMemoryToAccelerationStructureKHR = fn (     C.Device,     C.DeferredOperationKHR,     &CopyMemoryToAccelerationStructureInfoKHR) Result

pub fn copy_memory_to_acceleration_structure_khr(
    device                                          C.Device,
    deferred_operation                              C.DeferredOperationKHR,
    p_info                                          &CopyMemoryToAccelerationStructureInfoKHR) Result {
      f := VkCopyMemoryToAccelerationStructureKHR((*loader_p).get_sym('vkCopyMemoryToAccelerationStructureKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCopyMemoryToAccelerationStructureKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    deferred_operation,
    p_info)
}


type VkWriteAccelerationStructuresPropertiesKHR = fn (     C.Device,     u32,     &C.AccelerationStructureKHR,     QueryType,     usize,     voidptr,     usize) Result

pub fn write_acceleration_structures_properties_khr(
    device                                          C.Device,
    acceleration_structure_count                    u32,
    p_acceleration_structures                       &C.AccelerationStructureKHR,
    query_type                                      QueryType,
    data_size                                       usize,
    p_data                                          voidptr,
    stride                                          usize) Result {
      f := VkWriteAccelerationStructuresPropertiesKHR((*loader_p).get_sym('vkWriteAccelerationStructuresPropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkWriteAccelerationStructuresPropertiesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    acceleration_structure_count,
    p_acceleration_structures,
    query_type,
    data_size,
    p_data,
    stride)
}


type VkCmdCopyAccelerationStructureKHR = fn (     C.CommandBuffer,     &CopyAccelerationStructureInfoKHR) 

pub fn cmd_copy_acceleration_structure_khr(
    command_buffer                                  C.CommandBuffer,
    p_info                                          &CopyAccelerationStructureInfoKHR)  {
      f := VkCmdCopyAccelerationStructureKHR((*loader_p).get_sym('vkCmdCopyAccelerationStructureKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyAccelerationStructureKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_info)
}


type VkCmdCopyAccelerationStructureToMemoryKHR = fn (     C.CommandBuffer,     &CopyAccelerationStructureToMemoryInfoKHR) 

pub fn cmd_copy_acceleration_structure_to_memory_khr(
    command_buffer                                  C.CommandBuffer,
    p_info                                          &CopyAccelerationStructureToMemoryInfoKHR)  {
      f := VkCmdCopyAccelerationStructureToMemoryKHR((*loader_p).get_sym('vkCmdCopyAccelerationStructureToMemoryKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyAccelerationStructureToMemoryKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_info)
}


type VkCmdCopyMemoryToAccelerationStructureKHR = fn (     C.CommandBuffer,     &CopyMemoryToAccelerationStructureInfoKHR) 

pub fn cmd_copy_memory_to_acceleration_structure_khr(
    command_buffer                                  C.CommandBuffer,
    p_info                                          &CopyMemoryToAccelerationStructureInfoKHR)  {
      f := VkCmdCopyMemoryToAccelerationStructureKHR((*loader_p).get_sym('vkCmdCopyMemoryToAccelerationStructureKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdCopyMemoryToAccelerationStructureKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_info)
}


type VkGetAccelerationStructureDeviceAddressKHR = fn (     C.Device,     &AccelerationStructureDeviceAddressInfoKHR) DeviceAddress

pub fn get_acceleration_structure_device_address_khr(
    device                                          C.Device,
    p_info                                          &AccelerationStructureDeviceAddressInfoKHR) DeviceAddress {
      f := VkGetAccelerationStructureDeviceAddressKHR((*loader_p).get_sym("vkGetAccelerationStructureDeviceAddressKHR"
    ) or { 
        panic("Couldn't load symbol for 'vkGetAccelerationStructureDeviceAddressKHR': ${err}") })
    return f(
    device,
    p_info)
}


type VkCmdWriteAccelerationStructuresPropertiesKHR = fn (     C.CommandBuffer,     u32,     &C.AccelerationStructureKHR,     QueryType,     C.QueryPool,     u32) 

pub fn cmd_write_acceleration_structures_properties_khr(
    command_buffer                                  C.CommandBuffer,
    acceleration_structure_count                    u32,
    p_acceleration_structures                       &C.AccelerationStructureKHR,
    query_type                                      QueryType,
    query_pool                                      C.QueryPool,
    first_query                                     u32)  {
      f := VkCmdWriteAccelerationStructuresPropertiesKHR((*loader_p).get_sym('vkCmdWriteAccelerationStructuresPropertiesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdWriteAccelerationStructuresPropertiesKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    acceleration_structure_count,
    p_acceleration_structures,
    query_type,
    query_pool,
    first_query)
}


type VkGetDeviceAccelerationStructureCompatibilityKHR = fn (     C.Device,     &AccelerationStructureVersionInfoKHR,     &AccelerationStructureCompatibilityKHR) 

pub fn get_device_acceleration_structure_compatibility_khr(
    device                                          C.Device,
    p_version_info                                  &AccelerationStructureVersionInfoKHR,
    p_compatibility                                 &AccelerationStructureCompatibilityKHR)  {
      f := VkGetDeviceAccelerationStructureCompatibilityKHR((*loader_p).get_sym('vkGetDeviceAccelerationStructureCompatibilityKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetDeviceAccelerationStructureCompatibilityKHR': ${err}")
        return 
    })
    f(
    device,
    p_version_info,
    p_compatibility)
}


type VkGetAccelerationStructureBuildSizesKHR = fn (     C.Device,     AccelerationStructureBuildTypeKHR,     &AccelerationStructureBuildGeometryInfoKHR,     &u32,     &AccelerationStructureBuildSizesInfoKHR) 

pub fn get_acceleration_structure_build_sizes_khr(
    device                                          C.Device,
    build_type                                      AccelerationStructureBuildTypeKHR,
    p_build_info                                    &AccelerationStructureBuildGeometryInfoKHR,
    p_max_primitive_counts                          &u32,
    p_size_info                                     &AccelerationStructureBuildSizesInfoKHR)  {
      f := VkGetAccelerationStructureBuildSizesKHR((*loader_p).get_sym('vkGetAccelerationStructureBuildSizesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetAccelerationStructureBuildSizesKHR': ${err}")
        return 
    })
    f(
    device,
    build_type,
    p_build_info,
    p_max_primitive_counts,
    p_size_info)
}




// VK_KHR_ray_tracing_pipeline is a preprocessor guard. Do not pass it to API calls.
const khr_ray_tracing_pipeline = 1
pub const khr_ray_tracing_pipeline_spec_version = 1
pub const khr_ray_tracing_pipeline_extension_name = "VK_KHR_ray_tracing_pipeline"

pub enum ShaderGroupShaderKHR {
    shader_group_shader_general_khr = int(0)
    shader_group_shader_closest_hit_khr = int(1)
    shader_group_shader_any_hit_khr = int(2)
    shader_group_shader_intersection_khr = int(3)
    shader_group_shader_max_enum_khr = int(0x7FFFFFFF)
}

pub struct RayTracingShaderGroupCreateInfoKHR {
mut:
    s_type                                StructureType
    p_next                                voidptr
    vktype                                RayTracingShaderGroupTypeKHR
    general_shader                        u32
    closest_hit_shader                    u32
    any_hit_shader                        u32
    intersection_shader                   u32
    p_shader_group_capture_replay_handle  voidptr
} 

pub struct RayTracingPipelineInterfaceCreateInfoKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_pipeline_ray_payload_size u32
    max_pipeline_ray_hit_attribute_size u32
} 

pub struct RayTracingPipelineCreateInfoKHR {
mut:
    s_type                                                   StructureType
    p_next                                                   voidptr
    flags                                                    PipelineCreateFlags
    stage_count                                              u32
    p_stages                                                 &PipelineShaderStageCreateInfo
    group_count                                              u32
    p_groups                                                 &RayTracingShaderGroupCreateInfoKHR
    max_pipeline_ray_recursion_depth                         u32
    p_library_info                                           &PipelineLibraryCreateInfoKHR
    p_library_interface                                      &RayTracingPipelineInterfaceCreateInfoKHR
    p_dynamic_state                                          &PipelineDynamicStateCreateInfo
    layout                                                   C.PipelineLayout
    base_pipeline_handle                                     C.Pipeline
    base_pipeline_index                                      i32
} 

// PhysicalDeviceRayTracingPipelineFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRayTracingPipelineFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    ray_tracing_pipeline   Bool32
    ray_tracing_pipeline_shader_group_handle_capture_replay Bool32
    ray_tracing_pipeline_shader_group_handle_capture_replay_mixed Bool32
    ray_tracing_pipeline_trace_rays_indirect Bool32
    ray_traversal_primitive_culling Bool32
} 

// PhysicalDeviceRayTracingPipelinePropertiesKHR extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceRayTracingPipelinePropertiesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    shader_group_handle_size u32
    max_ray_recursion_depth u32
    max_shader_group_stride u32
    shader_group_base_alignment u32
    shader_group_handle_capture_replay_size u32
    max_ray_dispatch_invocation_count u32
    shader_group_handle_alignment u32
    max_ray_hit_attribute_size u32
} 

pub struct StridedDeviceAddressRegionKHR {
mut:
    device_address         DeviceAddress
    stride                 DeviceSize
    size                   DeviceSize
} 

pub struct TraceRaysIndirectCommandKHR {
mut:
    width           u32
    height          u32
    depth           u32
} 

type VkCmdTraceRaysKHR = fn (     C.CommandBuffer,     &StridedDeviceAddressRegionKHR,     &StridedDeviceAddressRegionKHR,     &StridedDeviceAddressRegionKHR,     &StridedDeviceAddressRegionKHR,     u32,     u32,     u32) 

pub fn cmd_trace_rays_khr(
    command_buffer                                  C.CommandBuffer,
    p_raygen_shader_binding_table                   &StridedDeviceAddressRegionKHR,
    p_miss_shader_binding_table                     &StridedDeviceAddressRegionKHR,
    p_hit_shader_binding_table                      &StridedDeviceAddressRegionKHR,
    p_callable_shader_binding_table                 &StridedDeviceAddressRegionKHR,
    width                                           u32,
    height                                          u32,
    depth                                           u32)  {
      f := VkCmdTraceRaysKHR((*loader_p).get_sym('vkCmdTraceRaysKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdTraceRaysKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_raygen_shader_binding_table,
    p_miss_shader_binding_table,
    p_hit_shader_binding_table,
    p_callable_shader_binding_table,
    width,
    height,
    depth)
}


type VkCreateRayTracingPipelinesKHR = fn (     C.Device,     C.DeferredOperationKHR,     C.PipelineCache,     u32,     &RayTracingPipelineCreateInfoKHR,     &AllocationCallbacks,     &C.Pipeline) Result

pub fn create_ray_tracing_pipelines_khr(
    device                                          C.Device,
    deferred_operation                              C.DeferredOperationKHR,
    pipeline_cache                                  C.PipelineCache,
    create_info_count                               u32,
    p_create_infos                                  &RayTracingPipelineCreateInfoKHR,
    p_allocator                                     &AllocationCallbacks,
    p_pipelines                                     &C.Pipeline) Result {
      f := VkCreateRayTracingPipelinesKHR((*loader_p).get_sym('vkCreateRayTracingPipelinesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCreateRayTracingPipelinesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    deferred_operation,
    pipeline_cache,
    create_info_count,
    p_create_infos,
    p_allocator,
    p_pipelines)
}


type VkGetRayTracingCaptureReplayShaderGroupHandlesKHR = fn (     C.Device,     C.Pipeline,     u32,     u32,     usize,     voidptr) Result

pub fn get_ray_tracing_capture_replay_shader_group_handles_khr(
    device                                          C.Device,
    pipeline                                        C.Pipeline,
    first_group                                     u32,
    group_count                                     u32,
    data_size                                       usize,
    p_data                                          voidptr) Result {
      f := VkGetRayTracingCaptureReplayShaderGroupHandlesKHR((*loader_p).get_sym('vkGetRayTracingCaptureReplayShaderGroupHandlesKHR'
    ) or { 
        println("Couldn't load symbol for 'vkGetRayTracingCaptureReplayShaderGroupHandlesKHR': ${err}")
        return Result.error_unknown
    })
    return f(
    device,
    pipeline,
    first_group,
    group_count,
    data_size,
    p_data)
}


type VkCmdTraceRaysIndirectKHR = fn (     C.CommandBuffer,     &StridedDeviceAddressRegionKHR,     &StridedDeviceAddressRegionKHR,     &StridedDeviceAddressRegionKHR,     &StridedDeviceAddressRegionKHR,     DeviceAddress) 

pub fn cmd_trace_rays_indirect_khr(
    command_buffer                                  C.CommandBuffer,
    p_raygen_shader_binding_table                   &StridedDeviceAddressRegionKHR,
    p_miss_shader_binding_table                     &StridedDeviceAddressRegionKHR,
    p_hit_shader_binding_table                      &StridedDeviceAddressRegionKHR,
    p_callable_shader_binding_table                 &StridedDeviceAddressRegionKHR,
    indirect_device_address                         DeviceAddress)  {
      f := VkCmdTraceRaysIndirectKHR((*loader_p).get_sym('vkCmdTraceRaysIndirectKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdTraceRaysIndirectKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    p_raygen_shader_binding_table,
    p_miss_shader_binding_table,
    p_hit_shader_binding_table,
    p_callable_shader_binding_table,
    indirect_device_address)
}


type VkGetRayTracingShaderGroupStackSizeKHR = fn (     C.Device,     C.Pipeline,     u32,     ShaderGroupShaderKHR) DeviceSize

pub fn get_ray_tracing_shader_group_stack_size_khr(
    device                                          C.Device,
    pipeline                                        C.Pipeline,
    group                                           u32,
    group_shader                                    ShaderGroupShaderKHR) DeviceSize {
      f := VkGetRayTracingShaderGroupStackSizeKHR((*loader_p).get_sym("vkGetRayTracingShaderGroupStackSizeKHR"
    ) or { 
        panic("Couldn't load symbol for 'vkGetRayTracingShaderGroupStackSizeKHR': ${err}") })
    return f(
    device,
    pipeline,
    group,
    group_shader)
}


type VkCmdSetRayTracingPipelineStackSizeKHR = fn (     C.CommandBuffer,     u32) 

pub fn cmd_set_ray_tracing_pipeline_stack_size_khr(
    command_buffer                                  C.CommandBuffer,
    pipeline_stack_size                             u32)  {
      f := VkCmdSetRayTracingPipelineStackSizeKHR((*loader_p).get_sym('vkCmdSetRayTracingPipelineStackSizeKHR'
    ) or { 
        println("Couldn't load symbol for 'vkCmdSetRayTracingPipelineStackSizeKHR': ${err}")
        return 
    })
    f(
    command_buffer,
    pipeline_stack_size)
}




// VK_KHR_ray_query is a preprocessor guard. Do not pass it to API calls.
const khr_ray_query = 1
pub const khr_ray_query_spec_version        = 1
pub const khr_ray_query_extension_name      = "VK_KHR_ray_query"
// PhysicalDeviceRayQueryFeaturesKHR extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceRayQueryFeaturesKHR {
mut:
    s_type                 StructureType
    p_next                 voidptr
    ray_query              Bool32
} 



// VK_EXT_mesh_shader is a preprocessor guard. Do not pass it to API calls.
const ext_mesh_shader = 1
pub const ext_mesh_shader_spec_version      = 1
pub const ext_mesh_shader_extension_name    = "VK_EXT_mesh_shader"
// PhysicalDeviceMeshShaderFeaturesEXT extends VkPhysicalDeviceFeatures2,VkDeviceCreateInfo
pub struct PhysicalDeviceMeshShaderFeaturesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    task_shader            Bool32
    mesh_shader            Bool32
    multiview_mesh_shader  Bool32
    primitive_fragment_shading_rate_mesh_shader Bool32
    mesh_shader_queries    Bool32
} 

// PhysicalDeviceMeshShaderPropertiesEXT extends VkPhysicalDeviceProperties2
pub struct PhysicalDeviceMeshShaderPropertiesEXT {
mut:
    s_type                 StructureType
    p_next                 voidptr
    max_task_work_group_total_count u32
    max_task_work_group_count []u32
    max_task_work_group_invocations u32
    max_task_work_group_size []u32
    max_task_payload_size  u32
    max_task_shared_memory_size u32
    max_task_payload_and_shared_memory_size u32
    max_mesh_work_group_total_count u32
    max_mesh_work_group_count []u32
    max_mesh_work_group_invocations u32
    max_mesh_work_group_size []u32
    max_mesh_shared_memory_size u32
    max_mesh_payload_and_shared_memory_size u32
    max_mesh_output_memory_size u32
    max_mesh_payload_and_output_memory_size u32
    max_mesh_output_components u32
    max_mesh_output_vertices u32
    max_mesh_output_primitives u32
    max_mesh_output_layers u32
    max_mesh_multiview_view_count u32
    mesh_output_per_vertex_granularity u32
    mesh_output_per_primitive_granularity u32
    max_preferred_task_work_group_invocations u32
    max_preferred_mesh_work_group_invocations u32
    prefers_local_invocation_vertex_output Bool32
    prefers_local_invocation_primitive_output Bool32
    prefers_compact_vertex_output Bool32
    prefers_compact_primitive_output Bool32
} 

pub struct DrawMeshTasksIndirectCommandEXT {
mut:
    group_count_x   u32
    group_count_y   u32
    group_count_z   u32
} 

type VkCmdDrawMeshTasksEXT = fn (     C.CommandBuffer,     u32,     u32,     u32) 

pub fn cmd_draw_mesh_tasks_ext(
    command_buffer                                  C.CommandBuffer,
    group_count_x                                   u32,
    group_count_y                                   u32,
    group_count_z                                   u32)  {
      f := VkCmdDrawMeshTasksEXT((*loader_p).get_sym('vkCmdDrawMeshTasksEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawMeshTasksEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    group_count_x,
    group_count_y,
    group_count_z)
}


type VkCmdDrawMeshTasksIndirectEXT = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_mesh_tasks_indirect_ext(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    draw_count                                      u32,
    stride                                          u32)  {
      f := VkCmdDrawMeshTasksIndirectEXT((*loader_p).get_sym('vkCmdDrawMeshTasksIndirectEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawMeshTasksIndirectEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    draw_count,
    stride)
}


type VkCmdDrawMeshTasksIndirectCountEXT = fn (     C.CommandBuffer,     C.Buffer,     DeviceSize,     C.Buffer,     DeviceSize,     u32,     u32) 

pub fn cmd_draw_mesh_tasks_indirect_count_ext(
    command_buffer                                  C.CommandBuffer,
    buffer                                          C.Buffer,
    offset                                          DeviceSize,
    count_buffer                                    C.Buffer,
    count_buffer_offset                             DeviceSize,
    max_draw_count                                  u32,
    stride                                          u32)  {
      f := VkCmdDrawMeshTasksIndirectCountEXT((*loader_p).get_sym('vkCmdDrawMeshTasksIndirectCountEXT'
    ) or { 
        println("Couldn't load symbol for 'vkCmdDrawMeshTasksIndirectCountEXT': ${err}")
        return 
    })
    f(
    command_buffer,
    buffer,
    offset,
    count_buffer,
    count_buffer_offset,
    max_draw_count,
    stride)
}


